-------------------------------------------------------------------------
-- Design unit: Memory
-- Description: Parametrizable memory
--      Synchronous read and write
-------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;
use work.Util_package.all;


entity VMemory is
    generic (
        DATA_WIDTH  : integer := 8;         -- Data bus width
        ADDR_WIDTH  : integer := 8;         -- Address bus width
        IMAGE       : string := "UNUSED"    -- Memory content to be loaded    (text file)
    );
    port (  
        clk         : in std_logic;
        we          : in std_logic;        -- Write Enable
        address     : in std_logic_vector (ADDR_WIDTH-1 downto 0);
        data_in     : in std_logic_vector (DATA_WIDTH-1 downto 0);
        data_out    : out std_logic_vector (DATA_WIDTH-1 downto 0)
    );
end VMemory;

architecture BLOCK_RAM of VMemory is
    
    type RamType is array (0 to (2**ADDR_WIDTH)-1) of std_logic_vector(DATA_WIDTH-1 downto 0);
    
    impure function InitRamFromFile (RamFileName : in string) return RamType is
        FILE RamFile : text is in RamFileName;
        variable RamFileLine : line;
        variable RAM : RamType;
        variable str : string(1 to 2);
    begin   
        for I in RamType'range loop
            readline (RamFile, RamFileLine);
            read (RamFileLine, str);
            RAM(I) := StringToStdLogicVector(str);
        end loop;
        return RAM;
    end function;
    
    signal RAM : RamType := InitRamFromFile(IMAGE);
   
    
    -- Teste resolução 640x480 (primeira e última colunas são brancas)
    --signal RAM : RamType := (
    --    -- 100 pixels (0-99) colunas vermelhas
    --    x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"A0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"A0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"A0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"A0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"A0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"A0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"A0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"A0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"A0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    --    
    --    -- 100 pixels (100-199) colunas verdes
    --    x"14",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"14",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"14",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"14",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"14",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"14",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"14",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"14",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"14",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"14",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    --
    --    -- 100 pixels (200-299) colunas vermelhas
    --    x"A0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"A0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"A0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"A0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"A0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"A0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"A0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"A0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"A0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"A0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    --    
    --    -- 100 pixels (300-399) colunas verdes
    --    x"14",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"14",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"14",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"14",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"14",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"14",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"14",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"14",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"14",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"14",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    --
    --    -- 100 pixels (400-499) colunas vermelhas
    --    x"A0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"A0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"A0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"A0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"A0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"A0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"A0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"A0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"A0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"A0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    --    
    --    -- 100 pixels (500-599) colunas verdes
    --    x"14",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"14",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"14",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"14",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"14",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"14",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"14",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"14",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"14",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"14",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    --
    --    -- 100 pixels (600-40) colunas vermelhas
    --    x"A0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"A0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"A0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"A0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF", x"03",
    --    
    --    others=>x"00");
        
    -- Teste resolução 800x600 (primeira e última colunas são brancas)    
    --signal RAM : RamType := (
    --    -- 100 pixels (0-99) colunas vermelhas
    --    x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"A0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"A0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"A0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"A0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"A0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"A0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"A0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"A0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"A0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    --    
    --    -- 100 pixels (100-199) colunas verdes
    --    x"14",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"14",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"14",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"14",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"14",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"14",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"14",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"14",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"14",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"14",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    --
    --    -- 100 pixels (200-299) colunas vermelhas
    --    x"A0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"A0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"A0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"A0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"A0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"A0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"A0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"A0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"A0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"A0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    --    
    --    -- 100 pixels (300-399) colunas verdes
    --    x"14",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"14",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"14",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"14",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"14",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"14",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"14",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"14",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"14",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"14",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    --
    --    -- 100 pixels (400-499) colunas vermelhas
    --    x"A0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"A0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"A0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"A0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"A0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"A0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"A0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"A0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"A0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"A0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    --    
    --    -- 100 pixels (500-599) colunas verdes
    --    x"14",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"14",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"14",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"14",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"14",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"14",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"14",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"14",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"14",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"14",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    --
    --    -- 100 pixels (600-699) colunas vermelhas
    --    x"A0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"A0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"A0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"A0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"A0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"A0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"A0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"A0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"A0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"A0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    --    
    --    -- 100 pixels (700-799) colunas verdes
    --    x"14",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"14",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"14",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"14",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"14",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"14",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"14",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"14",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"14",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", x"14",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",
    -- 
    --others=>x"00");
    
    -- surfer.bmp
--    signal RAM : RamType := (
--        x"09",x"09",x"EC",x"EC",x"EC",x"EC",x"EC",x"F4",x"F5",x"F5",x"F5",x"F5",x"09",x"09",x"09",x"F6",x"F6",x"09",x"09",x"09",x"09",x"07",x"09",x"09",x"F6",x"F6",x"F6",x"F6",x"F6",x"09",x"09",x"09",
--        x"09",x"09",x"09",x"09",x"EC",x"EC",x"EC",x"F4",x"EC",x"EC",x"EC",x"F5",x"F4",x"F5",x"09",x"A4",x"A4",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",
--        x"F5",x"09",x"09",x"09",x"F5",x"F5",x"F5",x"F5",x"F4",x"F4",x"F5",x"EC",x"EC",x"EC",x"92",x"41",x"00",x"A4",x"ED",x"F4",x"F4",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",
--        x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"F4",x"09",x"09",x"09",x"09",x"52",x"00",x"00",x"F7",x"ED",x"EC",x"E3",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"ED",x"09",x"09",x"09",x"09",
--        x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"F5",x"F5",x"F5",x"09",x"09",x"09",x"09",x"49",x"51",x"09",x"09",x"09",x"09",x"09",x"09",x"F4",x"EC",x"EC",x"E3",x"A3",x"E3",x"E3",x"E4",x"EC",
--        x"F5",x"F5",x"09",x"F5",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"EC",x"E4",x"EC",x"09",x"09",x"EC",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"F5",x"F5",x"EC",x"EC",x"EC",x"EC",
--        x"09",x"09",x"09",x"09",x"09",x"F5",x"F5",x"F5",x"F5",x"09",x"09",x"DA",x"91",x"91",x"89",x"EC",x"EC",x"EC",x"EB",x"EC",x"EC",x"F5",x"09",x"F4",x"F5",x"09",x"09",x"09",x"09",x"EC",x"EC",x"EC",
--        x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"F5",x"EC",x"E2",x"DA",x"91",x"40",x"40",x"DA",x"9B",x"F5",x"F4",x"EB",x"F4",x"EC",x"EC",x"EC",x"EC",x"09",x"09",x"09",x"09",x"F5",x"EC",x"EC",
--        x"F5",x"F5",x"09",x"09",x"09",x"09",x"F4",x"EC",x"ED",x"E3",x"DA",x"E3",x"91",x"48",x"00",x"49",x"EC",x"09",x"F4",x"09",x"07",x"F5",x"09",x"09",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"09",
--        x"F5",x"F5",x"ED",x"ED",x"F5",x"F5",x"EC",x"EC",x"EC",x"48",x"48",x"49",x"48",x"00",x"A3",x"92",x"92",x"EC",x"EB",x"A3",x"A3",x"E3",x"F4",x"EC",x"EC",x"EC",x"EC",x"EC",x"E3",x"E3",x"E3",x"E3",
--        x"F5",x"ED",x"EC",x"EC",x"EC",x"ED",x"ED",x"ED",x"ED",x"00",x"00",x"00",x"00",x"00",x"ED",x"09",x"89",x"9A",x"09",x"09",x"EC",x"E3",x"E3",x"EC",x"E3",x"E3",x"EC",x"EC",x"EC",x"EC",x"F5",x"F4",
--        x"09",x"09",x"F5",x"F5",x"ED",x"ED",x"EC",x"EC",x"ED",x"49",x"00",x"00",x"00",x"00",x"00",x"ED",x"09",x"92",x"A2",x"09",x"09",x"F5",x"09",x"09",x"EC",x"E4",x"EC",x"EC",x"E3",x"E3",x"EC",x"EC",
--        x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"ED",x"00",x"00",x"00",x"00",x"00",x"49",x"ED",x"F5",x"9B",x"4A",x"E5",x"07",x"ED",x"EC",x"F5",x"EC",x"ED",x"F5",x"EC",x"EC",x"EC",x"F5",
--        x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"F6",x"A4",x"00",x"00",x"52",x"00",x"00",x"49",x"F5",x"F5",x"52",x"52",x"EE",x"09",x"F5",x"F5",x"ED",x"EC",x"EC",x"EC",x"EC",x"ED",x"F5",
--        x"F6",x"F6",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"A3",x"00",x"9B",x"F6",x"F5",x"00",x"49",x"F5",x"09",x"07",x"ED",x"ED",x"F5",x"ED",x"ED",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",
--        x"FF",x"FF",x"F6",x"09",x"09",x"09",x"F5",x"F5",x"09",x"AC",x"00",x"52",x"F6",x"09",x"09",x"49",x"00",x"09",x"09",x"09",x"09",x"09",x"F5",x"09",x"F5",x"EC",x"ED",x"ED",x"ED",x"EC",x"ED",x"F5",
--        x"09",x"09",x"FF",x"FF",x"FF",x"F6",x"09",x"07",x"07",x"49",x"00",x"E4",x"09",x"09",x"09",x"51",x"00",x"ED",x"09",x"09",x"07",x"F5",x"09",x"09",x"09",x"09",x"09",x"09",x"F5",x"F5",x"EC",x"EC",
--        x"A3",x"E3",x"ED",x"09",x"F6",x"F6",x"F6",x"FF",x"ED",x"92",x"ED",x"ED",x"A3",x"E3",x"E3",x"9A",x"00",x"AC",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",
--        x"EC",x"E3",x"9B",x"A3",x"A3",x"E3",x"E3",x"E4",x"E4",x"EC",x"FF",x"FF",x"08",x"09",x"ED",x"9B",x"00",x"92",x"EC",x"EC",x"EC",x"EC",x"E3",x"EC",x"F5",x"F5",x"09",x"09",x"09",x"09",x"09",x"09",
--        x"09",x"09",x"ED",x"ED",x"EC",x"E3",x"9A",x"91",x"49",x"52",x"9C",x"F7",x"08",x"F6",x"FF",x"07",x"00",x"00",x"48",x"A3",x"EC",x"A3",x"DB",x"DA",x"E3",x"E3",x"EB",x"EB",x"EC",x"F5",x"F4",x"F5",
--        x"09",x"09",x"09",x"09",x"09",x"F5",x"F5",x"F5",x"51",x"00",x"49",x"52",x"92",x"9B",x"A4",x"A4",x"52",x"53",x"53",x"B7",x"BF",x"B7",x"08",x"07",x"07",x"F7",x"ED",x"F7",x"E4",x"E4",x"E3",x"E3",
--        x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"9A",x"40",x"91",x"EC",x"EC",x"E3",x"A3",x"00",x"49",x"52",x"A5",x"AF",x"6E",x"6F",x"B7",x"BF",x"B7",x"B7",x"BF",x"B7",x"07",x"F7",x"E3",x"E3",
--        x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"9A",x"48",x"A3",x"EC",x"F4",x"09",x"A3",x"00",x"E3",x"E4",x"E4",x"EC",x"A4",x"9B",x"9B",x"9A",x"E3",x"9B",x"9B",x"9B",x"DB",x"E3",x"E3",x"EC",
--        x"09",x"09",x"09",x"09",x"09",x"09",x"09",x"EC",x"92",x"49",x"A4",x"ED",x"F5",x"EC",x"51",x"52",x"F5",x"F5",x"09",x"09",x"09",x"07",x"09",x"F5",x"EC",x"EC",x"E4",x"EC",x"EC",x"EC",x"EC",x"E3",
--    others=>x"00");
    
    -- pam.bmp
--    signal RAM : RamType := (
--        x"5C",x"5C",x"5B",x"AC",x"F7",x"F4",x"F4",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"F4",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"F7",x"F7",x"F7",x"AC",x"A4",x"64",x"5C",x"5C",x"65",x"AE",x"A5",x"A5",x"A5",x"A5",x"AD",x"AD",x"A4",x"A4",x"64",x"5C",x"5B",x"53",x"53",x"53",x"53",x"53",x"53",x"53",x"53",x"13",x"53",x"53",x"53",x"53",x"53",x"53",x"53",x"53",x"53",x"52",x"52",x"52",x"52",x"52",x"0A",x"52",x"52",x"52",x"52",x"52",x"52",x"4A",x"4A",x"52", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", 
--        x"5C",x"5C",x"5B",x"A4",x"F7",x"EC",x"F4",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"F7",x"F7",x"F7",x"F7",x"F7",x"AC",x"A4",x"64",x"5C",x"5C",x"5C",x"65",x"AE",x"A6",x"AE",x"AE",x"AD",x"AD",x"A5",x"63",x"5B",x"5B",x"5B",x"5B",x"53",x"53",x"53",x"13",x"12",x"13",x"13",x"12",x"12",x"13",x"13",x"13",x"53",x"53",x"53",x"52",x"52",x"52",x"52",x"52",x"52",x"52",x"0A",x"0A",x"0A",x"0A",x"52",x"52",x"52",x"4A",x"52",x"52",x"4A", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"5C",x"5C",x"5B",x"A3",x"F7",x"EC",x"F4",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"F7",x"F7",x"F7",x"F7",x"F7",x"AD",x"A4",x"64",x"5C",x"5C",x"5C",x"5C",x"65",x"A5",x"65",x"A5",x"A5",x"A5",x"AD",x"AD",x"A5",x"A4",x"5B",x"5B",x"5B",x"5B",x"53",x"52",x"52",x"53",x"53",x"53",x"12",x"12",x"12",x"52",x"52",x"52",x"52",x"52",x"52",x"52",x"4A",x"0A",x"0A",x"0A",x"0A",x"0A",x"11",x"0A",x"0A",x"51",x"52",x"52",x"11",x"0A",x"52",x"0A", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"5C",x"5C",x"5C",x"5B",x"F7",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"F7",x"F7",x"AC",x"A4",x"A4",x"A4",x"5C",x"5C",x"5C",x"5C",x"64",x"65",x"65",x"5D",x"65",x"A5",x"A5",x"A5",x"AE",x"AE",x"AD",x"AD",x"AD",x"A4",x"A4",x"A4",x"5B",x"52",x"53",x"5B",x"52",x"52",x"52",x"52",x"52",x"52",x"52",x"52",x"4A",x"4A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"00",x"11",x"49",x"52",x"52",x"52",x"52",x"52",x"51",x"51",x"51",x"11", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"1C",x"5C",x"5C",x"5B",x"AC",x"F7",x"EC",x"F4",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"F7",x"F7",x"AC",x"A4",x"A4",x"5C",x"5C",x"5C",x"5C",x"5C",x"5C",x"65",x"5D",x"5C",x"5C",x"5C",x"65",x"A5",x"A6",x"AE",x"AE",x"AE",x"AE",x"AD",x"AD",x"AD",x"AD",x"A4",x"52",x"52",x"52",x"52",x"52",x"52",x"52",x"52",x"52",x"49",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"00",x"00",x"00",x"00",x"49",x"51",x"52",x"52",x"52",x"52",x"52",x"52",x"52",x"51",x"52", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"1D",x"5C",x"5C",x"5B",x"A4",x"F7",x"EC",x"F4",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"F7",x"AC",x"A4",x"64",x"5C",x"5C",x"5D",x"65",x"5C",x"5C",x"5C",x"5C",x"5C",x"5C",x"5C",x"5C",x"5C",x"5D",x"65",x"A5",x"AE",x"AE",x"B7",x"F7",x"AD",x"AD",x"A4",x"5B",x"52",x"49",x"51",x"52",x"52",x"52",x"5A",x"52",x"51",x"11",x"00",x"0A",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"0A",x"0A",x"52", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"1D",x"1C",x"5C",x"5C",x"A3",x"F7",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"F7",x"AC",x"A4",x"A4",x"5C",x"5C",x"5D",x"65",x"65",x"5D",x"5C",x"5D",x"5D",x"5C",x"5C",x"5C",x"5C",x"5C",x"5C",x"5C",x"5C",x"65",x"A6",x"AE",x"07",x"F7",x"F7",x"AD",x"A3",x"52",x"52",x"5A",x"5A",x"5A",x"5A",x"5A",x"52",x"51",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"48",x"48",x"48",x"49",x"49",x"49",x"49",x"49", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"1D",x"1D",x"5C",x"5C",x"5B",x"F7",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"AC",x"A4",x"A4",x"5C",x"5C",x"65",x"65",x"5D",x"65",x"5D",x"5D",x"65",x"65",x"5C",x"13",x"13",x"13",x"5C",x"5C",x"5C",x"5D",x"5D",x"65",x"A5",x"AE",x"F7",x"F7",x"AD",x"A4",x"5B",x"52",x"52",x"52",x"51",x"51",x"51",x"51",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"49",x"51",x"51", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"1D",x"1D",x"5C",x"5C",x"5B",x"AC",x"EC",x"EC",x"EC",x"EB",x"EB",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EB",x"EB",x"EC",x"EC",x"EC",x"EC",x"F7",x"A4",x"A4",x"64",x"5C",x"5D",x"66",x"66",x"66",x"5D",x"5C",x"65",x"65",x"5C",x"13",x"13",x"13",x"13",x"13",x"5C",x"5C",x"5D",x"AE",x"65",x"65",x"A5",x"AE",x"B6",x"AE",x"AD",x"5B",x"52",x"52",x"51",x"49",x"51",x"51",x"49",x"49",x"49",x"49",x"49",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"49",x"51",x"51",x"51",x"5A",x"5A",x"9A",x"A2",x"A2",x"A2",x"A3", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"1D",x"1D",x"5C",x"5C",x"5B",x"A4",x"ED",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"AC",x"AC",x"A4",x"5C",x"5C",x"5C",x"65",x"66",x"5D",x"5D",x"5C",x"5D",x"65",x"65",x"13",x"13",x"13",x"5B",x"5C",x"5C",x"5C",x"5C",x"53",x"65",x"B7",x"65",x"65",x"AE",x"AE",x"AE",x"AE",x"AD",x"A4",x"9B",x"52",x"51",x"49",x"49",x"48",x"49",x"51",x"49",x"51",x"51",x"51",x"51",x"5A",x"9A",x"9A",x"9A",x"A3",x"A3",x"A3",x"A3",x"A3",x"A3",x"A3",x"AB",x"A3",x"A2",x"AA",x"AA", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"1D",x"1C",x"5C",x"5C",x"5B",x"9C",x"F7",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"F7",x"F7",x"AC",x"AC",x"A4",x"5B",x"5C",x"5C",x"65",x"66",x"5D",x"14",x"5C",x"65",x"65",x"5C",x"13",x"13",x"13",x"13",x"65",x"65",x"65",x"65",x"5C",x"5D",x"B7",x"65",x"65",x"AE",x"AE",x"AE",x"B6",x"B6",x"AD",x"A4",x"A3",x"5B",x"5A",x"5A",x"5A",x"9A",x"A3",x"9A",x"A3",x"A3",x"A3",x"A3",x"A3",x"A3",x"A3",x"AB",x"AB",x"AB",x"A3",x"A3",x"A3",x"A3",x"A3",x"A3",x"EB",x"EB",x"EB",x"EA", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"1D",x"1C",x"5C",x"5C",x"5C",x"5B",x"A4",x"A4",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"F7",x"F7",x"F7",x"AD",x"A4",x"5B",x"5B",x"5C",x"65",x"65",x"5D",x"5C",x"5D",x"5D",x"66",x"65",x"5C",x"5C",x"5C",x"54",x"14",x"5C",x"AE",x"AE",x"AE",x"65",x"5D",x"AE",x"65",x"65",x"AE",x"AF",x"AE",x"AE",x"B6",x"F7",x"AD",x"AC",x"A4",x"A3",x"AC",x"AC",x"AC",x"EC",x"AC",x"AB",x"EB",x"EB",x"EB",x"EB",x"AB",x"AB",x"AB",x"A3",x"A3",x"A3",x"A3",x"A3",x"A3",x"A3",x"A3",x"A3",x"E2",x"E3",x"E2", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"1C",x"1C",x"5C",x"5C",x"5C",x"5B",x"5B",x"9B",x"A4",x"AC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"F7",x"F7",x"AD",x"A4",x"5C",x"53",x"5C",x"65",x"65",x"5D",x"5D",x"5C",x"5D",x"66",x"AE",x"5D",x"5D",x"66",x"65",x"5D",x"5D",x"5C",x"66",x"AE",x"AF",x"AE",x"65",x"AE",x"AE",x"5D",x"66",x"AF",x"AE",x"AE",x"B6",x"F7",x"F7",x"AC",x"AC",x"AC",x"EC",x"AC",x"AB",x"AB",x"AB",x"AB",x"AB",x"AB",x"AB",x"AB",x"AB",x"AB",x"A3",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"A3",x"E3",x"E3",x"EB", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"1C",x"1C",x"5C",x"5C",x"5C",x"5C",x"53",x"5B",x"5B",x"A3",x"A3",x"AC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"F7",x"F7",x"A5",x"5C",x"5C",x"5C",x"5D",x"66",x"65",x"5D",x"5D",x"5D",x"5D",x"66",x"AF",x"5D",x"5D",x"66",x"5D",x"5D",x"5D",x"5D",x"5C",x"A6",x"B7",x"AE",x"AE",x"AE",x"AE",x"5D",x"66",x"AF",x"AF",x"AE",x"AE",x"07",x"F7",x"F7",x"AC",x"EC",x"EC",x"AB",x"AB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"E3",x"EB",x"E3",x"E3",x"E3",x"E3",x"EB",x"EB", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"1C",x"5D",x"5C",x"5C",x"5C",x"5C",x"5B",x"5B",x"5A",x"5A",x"5A",x"A3",x"A3",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"F7",x"AD",x"A4",x"5C",x"5C",x"5C",x"65",x"AE",x"66",x"5D",x"5D",x"5D",x"65",x"A6",x"AF",x"66",x"5E",x"66",x"5E",x"66",x"5E",x"5E",x"55",x"66",x"AF",x"B7",x"AF",x"AE",x"AE",x"66",x"66",x"AF",x"B7",x"AE",x"AE",x"07",x"F7",x"F7",x"EC",x"EC",x"EC",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"E3",x"EB",x"EB",x"EB",x"EA",x"AA", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"1C",x"5D",x"5C",x"5C",x"5C",x"5C",x"5C",x"A4",x"5B",x"5A",x"5A",x"5A",x"9A",x"A3",x"A4",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"F7",x"AD",x"64",x"5C",x"5C",x"5C",x"66",x"AF",x"66",x"5C",x"5C",x"5D",x"66",x"AF",x"AF",x"5E",x"5E",x"66",x"66",x"A7",x"66",x"66",x"5E",x"54",x"A6",x"B7",x"AF",x"AE",x"B7",x"66",x"66",x"AF",x"B7",x"AE",x"AE",x"07",x"07",x"F7",x"AC",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EA",x"EA",x"AA", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"1C",x"5D",x"1C",x"5C",x"5D",x"5C",x"5C",x"AD",x"AC",x"A3",x"A3",x"9A",x"5A",x"5A",x"9B",x"A3",x"AB",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"F7",x"F7",x"A5",x"65",x"65",x"54",x"5C",x"A6",x"AE",x"65",x"5D",x"65",x"5C",x"A6",x"AF",x"A7",x"66",x"66",x"66",x"66",x"AF",x"A7",x"A7",x"66",x"5D",x"65",x"B7",x"B7",x"AE",x"B7",x"AE",x"AF",x"AF",x"B7",x"B7",x"AE",x"B6",x"F7",x"F7",x"F7",x"EC",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"E2",x"A2",x"E2",x"EA", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"1C",x"5D",x"1C",x"5C",x"5D",x"5C",x"5C",x"AD",x"F7",x"AC",x"AC",x"A3",x"A3",x"9A",x"5A",x"5A",x"9A",x"A3",x"AC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"F7",x"F7",x"A5",x"5D",x"5D",x"54",x"5D",x"AE",x"AE",x"A6",x"5D",x"65",x"5D",x"AF",x"AF",x"66",x"5E",x"66",x"66",x"66",x"AF",x"A7",x"A7",x"66",x"5D",x"5D",x"AF",x"B7",x"AE",x"AF",x"A6",x"AE",x"AF",x"B7",x"B7",x"AE",x"AE",x"07",x"F7",x"F7",x"EC",x"EC",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"A2",x"A2",x"A2",x"E2", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"1C",x"5D",x"1C",x"5C",x"5D",x"5C",x"5C",x"A4",x"F7",x"F7",x"EC",x"EC",x"AC",x"A3",x"9B",x"5A",x"5A",x"5A",x"9A",x"A3",x"AC",x"F7",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"F7",x"AD",x"A5",x"5C",x"5D",x"5C",x"65",x"AF",x"AE",x"AE",x"5D",x"5D",x"65",x"AF",x"AF",x"66",x"5D",x"66",x"66",x"66",x"A7",x"A7",x"A7",x"66",x"5D",x"5D",x"AF",x"B7",x"AE",x"AF",x"A6",x"65",x"AF",x"B7",x"B7",x"AE",x"AD",x"07",x"F7",x"F7",x"EC",x"EC",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"A2",x"A2",x"A2",x"E2", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"1C",x"5D",x"1C",x"5C",x"5C",x"5C",x"5C",x"A4",x"AC",x"F7",x"EC",x"EC",x"EC",x"F7",x"AC",x"A4",x"A3",x"5A",x"5A",x"5A",x"A3",x"A3",x"AC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"F7",x"AC",x"A5",x"A4",x"5C",x"5D",x"5C",x"A6",x"AF",x"AE",x"A6",x"5D",x"5D",x"AE",x"A6",x"AE",x"66",x"66",x"66",x"66",x"66",x"AF",x"A7",x"AF",x"A7",x"66",x"5D",x"A6",x"B7",x"AF",x"AF",x"AE",x"5D",x"AE",x"AF",x"B7",x"B7",x"AD",x"07",x"F7",x"F7",x"F7",x"EC",x"EC",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"E2",x"E2",x"E2",x"EB", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"1C",x"1C",x"5C",x"5D",x"5C",x"5C",x"5C",x"5B",x"AC",x"F7",x"EC",x"EC",x"EC",x"EC",x"F7",x"F7",x"AC",x"A3",x"9B",x"5A",x"5A",x"5A",x"A3",x"A3",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"F7",x"A4",x"A4",x"A5",x"5C",x"5D",x"5D",x"AE",x"AF",x"AF",x"65",x"5D",x"5D",x"AF",x"66",x"66",x"66",x"66",x"66",x"66",x"A7",x"AF",x"AF",x"AF",x"AF",x"66",x"5D",x"65",x"AE",x"AE",x"AE",x"AF",x"65",x"AF",x"AE",x"AF",x"B7",x"AD",x"07",x"F7",x"F7",x"F7",x"EC",x"EC",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"5D",x"1C",x"5D",x"5D",x"5C",x"5C",x"5C",x"5B",x"AC",x"F7",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"F7",x"AC",x"A4",x"A3",x"9B",x"5A",x"5A",x"5A",x"A3",x"A3",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"F7",x"A4",x"A4",x"A5",x"5D",x"5D",x"5D",x"AF",x"AE",x"AE",x"5C",x"65",x"65",x"AF",x"5D",x"66",x"65",x"65",x"5D",x"5D",x"66",x"66",x"AF",x"A6",x"A6",x"66",x"5C",x"5D",x"A6",x"AE",x"AE",x"AF",x"66",x"AF",x"AF",x"AE",x"B7",x"AE",x"07",x"07",x"F7",x"F7",x"F7",x"EC",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"5D",x"1C",x"5C",x"5D",x"5C",x"5C",x"5C",x"5B",x"A4",x"AC",x"F4",x"EC",x"EC",x"EC",x"EC",x"EC",x"F7",x"F7",x"F7",x"AC",x"AC",x"A3",x"9A",x"5A",x"9A",x"9A",x"A3",x"A3",x"EC",x"EC",x"EC",x"EC",x"AC",x"F7",x"A4",x"A4",x"A5",x"5D",x"5D",x"65",x"B7",x"AE",x"A6",x"5D",x"65",x"AE",x"66",x"5D",x"65",x"5C",x"5D",x"5D",x"5C",x"5D",x"5D",x"66",x"A6",x"66",x"5D",x"14",x"14",x"66",x"A6",x"AE",x"66",x"66",x"AF",x"AF",x"AF",x"AF",x"AE",x"B6",x"B6",x"F7",x"F7",x"F7",x"EC",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"5D",x"1C",x"5C",x"5D",x"5C",x"5C",x"5C",x"5B",x"A4",x"F7",x"F4",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"F7",x"EC",x"EC",x"AB",x"A3",x"9A",x"9A",x"5A",x"9A",x"A3",x"AC",x"AC",x"AC",x"F7",x"F7",x"A4",x"64",x"A5",x"5D",x"5D",x"5D",x"B7",x"A6",x"65",x"65",x"65",x"AF",x"66",x"5D",x"14",x"0B",x"14",x"5D",x"5D",x"54",x"54",x"66",x"AF",x"66",x"5D",x"0B",x"14",x"5D",x"66",x"66",x"66",x"5D",x"A6",x"AF",x"AF",x"AE",x"A5",x"AE",x"B6",x"07",x"F7",x"F7",x"AC",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"A2",x"E2",x"E2",x"EA", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"5C",x"5C",x"1C",x"5C",x"5C",x"5C",x"5C",x"5B",x"A3",x"F5",x"EC",x"F4",x"EB",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"AB",x"A3",x"9A",x"5A",x"5A",x"5A",x"A3",x"A4",x"AD",x"AD",x"A5",x"A5",x"5C",x"5D",x"5D",x"66",x"AF",x"66",x"A6",x"5D",x"A6",x"A6",x"66",x"66",x"54",x"54",x"5C",x"66",x"66",x"5D",x"5D",x"66",x"AF",x"66",x"5D",x"54",x"54",x"5D",x"66",x"66",x"66",x"66",x"66",x"AE",x"AF",x"B7",x"AE",x"AE",x"AE",x"AE",x"07",x"AC",x"F7",x"AB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"E2",x"E2",x"EA",x"EA", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"5C",x"5C",x"1C",x"5C",x"5C",x"5C",x"5C",x"5B",x"5B",x"F7",x"EC",x"F4",x"EB",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"F7",x"AC",x"A4",x"A3",x"5A",x"5A",x"5A",x"5B",x"A4",x"A4",x"A5",x"A5",x"5C",x"5D",x"5D",x"AE",x"AE",x"A6",x"AE",x"65",x"66",x"66",x"A6",x"5D",x"5D",x"65",x"66",x"66",x"A6",x"5D",x"5D",x"5D",x"AF",x"AF",x"66",x"66",x"66",x"66",x"66",x"66",x"5E",x"66",x"66",x"66",x"AE",x"AF",x"AE",x"AE",x"AE",x"AE",x"07",x"F7",x"AC",x"AB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EA",x"EA",x"EA",x"EA", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"5C",x"5C",x"1C",x"1C",x"5C",x"5C",x"5C",x"5B",x"5B",x"AC",x"EC",x"F4",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"F7",x"F7",x"AC",x"A4",x"9B",x"5B",x"5B",x"5C",x"64",x"65",x"A5",x"5C",x"5D",x"65",x"AF",x"AE",x"AE",x"AE",x"AE",x"66",x"66",x"AF",x"5D",x"66",x"A6",x"A6",x"A7",x"66",x"66",x"5D",x"5D",x"AF",x"AF",x"AF",x"AF",x"A7",x"A7",x"66",x"66",x"5E",x"66",x"66",x"66",x"66",x"AE",x"AE",x"AE",x"AE",x"AE",x"AE",x"F7",x"AC",x"EC",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EA",x"EA",x"EA", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"5C",x"5C",x"1C",x"1C",x"1C",x"5C",x"5C",x"5B",x"5B",x"A4",x"F7",x"F4",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"F7",x"F7",x"F7",x"F7",x"AC",x"A4",x"A3",x"5C",x"64",x"65",x"65",x"5C",x"5D",x"66",x"AE",x"AF",x"AE",x"A6",x"A6",x"65",x"66",x"AF",x"66",x"5E",x"66",x"A7",x"A7",x"66",x"5E",x"5D",x"66",x"A7",x"AF",x"AF",x"AF",x"AF",x"AF",x"A7",x"66",x"66",x"5D",x"66",x"66",x"66",x"66",x"66",x"AF",x"AE",x"AE",x"AE",x"F7",x"AC",x"EC",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"5C",x"5C",x"5C",x"1C",x"14",x"5C",x"5C",x"5B",x"5B",x"A3",x"F7",x"F4",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"ED",x"F7",x"F7",x"A4",x"A4",x"A5",x"65",x"5D",x"5D",x"65",x"66",x"66",x"AF",x"AE",x"AE",x"65",x"65",x"66",x"66",x"A7",x"5E",x"66",x"67",x"A7",x"66",x"5D",x"5D",x"66",x"AF",x"AF",x"AF",x"A7",x"AF",x"AF",x"A7",x"66",x"66",x"15",x"5D",x"66",x"A6",x"A6",x"65",x"A6",x"AE",x"AE",x"AE",x"AE",x"AD",x"F7",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EA",x"EA",x"EA",x"EA", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"5C",x"5C",x"5C",x"1C",x"14",x"5C",x"5C",x"5B",x"5B",x"5B",x"F7",x"F4",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"F7",x"A4",x"A5",x"65",x"5D",x"5D",x"66",x"66",x"66",x"AF",x"AE",x"AE",x"65",x"65",x"66",x"5D",x"66",x"5E",x"5E",x"67",x"67",x"5E",x"15",x"15",x"5E",x"67",x"67",x"67",x"67",x"AF",x"AF",x"67",x"66",x"5D",x"15",x"5D",x"66",x"A6",x"AE",x"AE",x"65",x"A6",x"AE",x"AE",x"AE",x"F7",x"AC",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"E3",x"E3",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"5C",x"5C",x"5C",x"1C",x"1C",x"5C",x"5C",x"5B",x"5B",x"5B",x"AC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"F7",x"A4",x"A6",x"65",x"65",x"66",x"66",x"5D",x"66",x"AF",x"AF",x"AE",x"65",x"65",x"66",x"5D",x"5D",x"5D",x"5E",x"5E",x"5E",x"5E",x"55",x"55",x"5E",x"66",x"67",x"67",x"67",x"67",x"67",x"67",x"66",x"5D",x"5D",x"66",x"66",x"A6",x"AE",x"AE",x"65",x"66",x"A6",x"AE",x"AE",x"F7",x"AC",x"A3",x"A3",x"E3",x"A3",x"A3",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"5C",x"5C",x"5C",x"1C",x"1C",x"1C",x"5C",x"5C",x"5B",x"5A",x"AC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"AC",x"A4",x"AE",x"65",x"A6",x"AF",x"66",x"5D",x"AE",x"AF",x"AF",x"A6",x"66",x"5D",x"66",x"A6",x"15",x"55",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"66",x"67",x"AF",x"AF",x"67",x"67",x"66",x"66",x"5D",x"1D",x"66",x"AE",x"66",x"AE",x"66",x"65",x"66",x"66",x"AE",x"AE",x"F7",x"A4",x"A3",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"5C",x"5C",x"5C",x"1C",x"1C",x"1C",x"5C",x"5C",x"5B",x"5B",x"A3",x"F7",x"EC",x"EB",x"EC",x"F4",x"F4",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EC",x"AC",x"A5",x"65",x"66",x"AE",x"66",x"66",x"66",x"AE",x"AF",x"AF",x"65",x"66",x"5C",x"5D",x"A6",x"5D",x"55",x"5D",x"5E",x"5D",x"55",x"55",x"5D",x"5E",x"5E",x"66",x"66",x"A7",x"67",x"5E",x"66",x"66",x"5D",x"5D",x"66",x"AF",x"66",x"66",x"66",x"5D",x"65",x"65",x"AE",x"AE",x"AE",x"A4",x"9B",x"9B",x"9A",x"A2",x"A2",x"A2",x"A2",x"9A",x"9A",x"9A",x"9A",x"A2",x"A2",x"A2",x"99",x"A2",x"99",x"A2",x"A2",x"A2",x"A2",x"A2", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"5C",x"5C",x"5C",x"1C",x"1C",x"1C",x"1C",x"5C",x"5B",x"5B",x"A3",x"AC",x"AB",x"AB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EB",x"EA",x"EA",x"EA",x"EA",x"E3",x"A3",x"A3",x"A4",x"A5",x"65",x"66",x"66",x"66",x"66",x"66",x"AF",x"B7",x"AE",x"A6",x"5D",x"54",x"5D",x"A6",x"5D",x"55",x"5D",x"5E",x"5D",x"55",x"15",x"5D",x"66",x"5E",x"5E",x"5D",x"5E",x"66",x"5E",x"66",x"5E",x"5D",x"5D",x"66",x"AF",x"66",x"66",x"66",x"65",x"65",x"65",x"AE",x"AE",x"AE",x"A4",x"64",x"A4",x"A3",x"A3",x"5A",x"52",x"52",x"52",x"52",x"5A",x"A3",x"A3",x"A2",x"A3",x"A2",x"A3",x"9A",x"A3",x"A2",x"A2",x"A2",x"A2", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"5C",x"5C",x"5C",x"5C",x"1C",x"1C",x"1C",x"5C",x"5C",x"5B",x"5B",x"A3",x"A3",x"A2",x"A2",x"A2",x"EB",x"E3",x"A2",x"A2",x"A3",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A3",x"A3",x"A4",x"AD",x"65",x"65",x"65",x"66",x"66",x"AE",x"AF",x"B7",x"AE",x"AE",x"5C",x"5D",x"5D",x"66",x"5E",x"54",x"5D",x"5D",x"5D",x"55",x"15",x"5D",x"66",x"66",x"5E",x"5E",x"5E",x"A7",x"A7",x"A6",x"5D",x"55",x"5D",x"66",x"66",x"66",x"66",x"66",x"66",x"65",x"65",x"AE",x"AE",x"AE",x"A5",x"5C",x"9C",x"5C",x"54",x"53",x"53",x"53",x"4A",x"4A",x"52",x"F7",x"ED",x"A4",x"9B",x"5B",x"A4",x"9C",x"9C",x"A4",x"9C",x"9C",x"9C", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"5C",x"5C",x"5C",x"5C",x"1C",x"1C",x"1C",x"5C",x"5C",x"5B",x"5B",x"A3",x"A3",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A3",x"A3",x"A4",x"AD",x"AE",x"65",x"65",x"65",x"66",x"66",x"A6",x"AF",x"AF",x"AF",x"66",x"5C",x"5D",x"5D",x"5D",x"66",x"55",x"5D",x"5D",x"5D",x"5D",x"5D",x"5D",x"5E",x"5E",x"5E",x"66",x"A7",x"A7",x"66",x"5E",x"55",x"55",x"5D",x"66",x"66",x"5D",x"5D",x"66",x"66",x"A6",x"AE",x"AF",x"AE",x"AF",x"5C",x"54",x"53",x"4C",x"4C",x"4C",x"54",x"5D",x"54",x"53",x"52",x"53",x"F7",x"07",x"F7",x"5C",x"53",x"54",x"55",x"5C",x"54",x"53",x"54", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"5C",x"5C",x"5C",x"5C",x"1C",x"1C",x"5C",x"5C",x"5C",x"5B",x"5B",x"9B",x"A3",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A3",x"A3",x"A3",x"AD",x"AE",x"65",x"65",x"5D",x"65",x"66",x"66",x"A6",x"AF",x"AE",x"AF",x"65",x"5D",x"5D",x"5D",x"5E",x"5E",x"14",x"15",x"5D",x"5D",x"5E",x"5E",x"5E",x"5E",x"66",x"66",x"A7",x"AF",x"A6",x"5D",x"14",x"14",x"5D",x"5E",x"66",x"5E",x"5D",x"5E",x"66",x"66",x"66",x"AE",x"AF",x"AF",x"AF",x"5D",x"54",x"4C",x"0C",x"0C",x"0C",x"55",x"5D",x"54",x"53",x"5B",x"52",x"5B",x"AD",x"07",x"AE",x"54",x"4C",x"9E",x"54",x"4C",x"0B",x"0B", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"5C",x"5C",x"5C",x"5C",x"1C",x"5C",x"5C",x"5C",x"5C",x"5B",x"5B",x"5B",x"A3",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A3",x"A3",x"A4",x"AD",x"AE",x"5D",x"5D",x"5D",x"66",x"66",x"66",x"66",x"AF",x"AF",x"AE",x"5D",x"66",x"14",x"5D",x"66",x"5D",x"14",x"14",x"15",x"5D",x"5D",x"5E",x"66",x"67",x"AF",x"A7",x"AF",x"A7",x"5E",x"54",x"14",x"14",x"5E",x"5E",x"5E",x"5D",x"5D",x"66",x"66",x"6F",x"66",x"66",x"AF",x"A6",x"AF",x"55",x"54",x"55",x"0D",x"0C",x"0C",x"0C",x"54",x"54",x"53",x"53",x"5B",x"12",x"12",x"64",x"B7",x"A6",x"5D",x"5D",x"55",x"54",x"0B",x"0B", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"5C",x"5C",x"5C",x"14",x"14",x"5C",x"5C",x"5C",x"5C",x"5C",x"5B",x"5B",x"A3",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A3",x"A3",x"A4",x"AD",x"AD",x"A5",x"65",x"5D",x"5D",x"66",x"66",x"66",x"66",x"A7",x"A6",x"66",x"65",x"65",x"5D",x"66",x"66",x"14",x"14",x"15",x"15",x"15",x"15",x"5E",x"5E",x"67",x"A7",x"66",x"67",x"5E",x"54",x"14",x"0B",x"14",x"5E",x"5E",x"5D",x"5D",x"66",x"66",x"66",x"6E",x"AE",x"AF",x"AF",x"66",x"A7",x"4C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"54",x"13",x"0A",x"52",x"0A",x"0A",x"0A",x"52",x"A5",x"5C",x"53",x"13",x"54",x"53",x"13",x"0B", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"5C",x"5C",x"1C",x"14",x"14",x"5C",x"5C",x"5C",x"5C",x"5C",x"5B",x"5B",x"A3",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A3",x"A3",x"A3",x"A4",x"AD",x"A5",x"5D",x"66",x"66",x"66",x"5E",x"5E",x"66",x"66",x"A7",x"5D",x"AE",x"66",x"5D",x"AF",x"AF",x"5D",x"55",x"5D",x"15",x"15",x"15",x"55",x"5E",x"5E",x"5E",x"5E",x"66",x"A7",x"5D",x"14",x"14",x"14",x"54",x"5D",x"5D",x"5D",x"5D",x"66",x"6E",x"66",x"66",x"66",x"AE",x"AF",x"5E",x"A7",x"0C",x"0C",x"4C",x"0B",x"0C",x"0B",x"0B",x"0B",x"0B",x"0A",x"52",x"0A",x"0A",x"0A",x"0A",x"5B",x"53",x"0A",x"13",x"0B",x"13",x"13",x"13", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"5C",x"5C",x"5C",x"5C",x"54",x"54",x"5C",x"5C",x"5C",x"5C",x"5B",x"5B",x"A3",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A3",x"A3",x"AC",x"AD",x"65",x"65",x"66",x"66",x"5E",x"5E",x"5D",x"66",x"66",x"5E",x"AF",x"66",x"66",x"66",x"66",x"66",x"5D",x"5D",x"55",x"5D",x"5E",x"5D",x"15",x"5E",x"5E",x"66",x"67",x"67",x"67",x"67",x"5D",x"14",x"14",x"54",x"5D",x"5D",x"5D",x"5D",x"66",x"66",x"66",x"AE",x"66",x"66",x"AF",x"AE",x"AF",x"A6",x"0C",x"0C",x"0C",x"0B",x"0C",x"0C",x"0B",x"0B",x"4B",x"0B",x"0A",x"0A",x"0A",x"0A",x"0A",x"12",x"0B",x"0A",x"0B",x"0B",x"0B",x"0B",x"0B", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"5C",x"5C",x"5C",x"5C",x"54",x"54",x"5C",x"5C",x"5C",x"5C",x"5B",x"5B",x"A3",x"A3",x"A2",x"A2",x"A2",x"A2",x"A2",x"A1",x"A1",x"A1",x"A2",x"A2",x"A3",x"A3",x"A4",x"A5",x"65",x"5C",x"66",x"66",x"AF",x"5E",x"5D",x"5D",x"66",x"67",x"66",x"A7",x"5D",x"66",x"66",x"66",x"66",x"5D",x"5D",x"5D",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"67",x"67",x"67",x"67",x"5E",x"14",x"14",x"54",x"5D",x"5D",x"5D",x"66",x"6E",x"66",x"65",x"6E",x"66",x"66",x"AF",x"AF",x"AF",x"A6",x"0C",x"0C",x"0C",x"0C",x"0C",x"0B",x"0B",x"4B",x"4B",x"4B",x"4A",x"0A",x"0A",x"0A",x"0A",x"4B",x"4B",x"4B",x"4B",x"0B",x"0B",x"0B",x"0B", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"1C",x"5C",x"5C",x"5C",x"5C",x"5C",x"5C",x"5C",x"5C",x"5C",x"5B",x"5B",x"9B",x"A3",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A3",x"A4",x"A4",x"A5",x"65",x"65",x"66",x"66",x"66",x"5D",x"5D",x"5D",x"5E",x"5E",x"5E",x"67",x"5D",x"66",x"AF",x"66",x"5E",x"5D",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"66",x"5D",x"14",x"54",x"5D",x"5D",x"66",x"66",x"6E",x"66",x"66",x"AE",x"66",x"66",x"AF",x"AF",x"AF",x"A6",x"14",x"0B",x"0C",x"4C",x"4C",x"4C",x"4B",x"54",x"54",x"53",x"4A",x"0A",x"0A",x"0A",x"0A",x"4B",x"0B",x"0B",x"0B",x"53",x"53",x"4B",x"0B", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"14",x"1C",x"5C",x"5C",x"5C",x"5C",x"5C",x"5C",x"5C",x"5C",x"5C",x"5B",x"5B",x"A3",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A3",x"A4",x"64",x"65",x"66",x"AF",x"66",x"5D",x"66",x"5D",x"5D",x"5D",x"5E",x"5E",x"5E",x"67",x"5E",x"66",x"66",x"5E",x"5D",x"5D",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"67",x"67",x"67",x"67",x"67",x"67",x"66",x"5D",x"14",x"14",x"5D",x"5D",x"5D",x"66",x"AF",x"AF",x"AF",x"AE",x"66",x"66",x"AE",x"AE",x"AE",x"A6",x"14",x"0B",x"0B",x"0B",x"4C",x"4B",x"4B",x"53",x"53",x"4A",x"0A",x"49",x"49",x"52",x"52",x"4B",x"4B",x"4B",x"4B",x"53",x"53",x"4B",x"4B", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"14",x"14",x"5C",x"5C",x"5B",x"53",x"54",x"5C",x"5C",x"5C",x"5C",x"5B",x"5B",x"A3",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A3",x"9B",x"AD",x"65",x"65",x"AE",x"AF",x"5D",x"5D",x"66",x"5D",x"15",x"5D",x"5E",x"5E",x"66",x"66",x"66",x"66",x"66",x"5E",x"5D",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"5E",x"15",x"15",x"5D",x"5D",x"5D",x"66",x"AF",x"B7",x"AF",x"66",x"5D",x"66",x"66",x"A6",x"A6",x"A6",x"5C",x"13",x"0B",x"0B",x"4B",x"0B",x"0B",x"53",x"52",x"0A",x"0A",x"11",x"11",x"12",x"0A",x"0A",x"0B",x"0B",x"0B",x"0A",x"0A",x"0A",x"0A", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"14",x"14",x"54",x"54",x"53",x"53",x"53",x"54",x"14",x"5C",x"5C",x"5B",x"5B",x"A3",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A3",x"A3",x"A4",x"AE",x"A6",x"5D",x"AF",x"AF",x"5D",x"66",x"66",x"5D",x"5D",x"66",x"5E",x"5E",x"67",x"66",x"66",x"67",x"66",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"67",x"67",x"67",x"5F",x"5F",x"67",x"67",x"67",x"67",x"5E",x"5D",x"15",x"5D",x"54",x"5D",x"AF",x"AF",x"AF",x"67",x"5D",x"66",x"66",x"66",x"66",x"66",x"AE",x"5D",x"5C",x"54",x"5C",x"54",x"53",x"0A",x"0A",x"0A",x"0A",x"0A",x"52",x"52",x"53",x"53",x"53",x"13",x"13",x"13",x"53",x"53",x"53",x"5B", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"14",x"14",x"54",x"53",x"53",x"53",x"53",x"54",x"14",x"5C",x"5C",x"5B",x"5B",x"A3",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A3",x"A3",x"A4",x"A5",x"A6",x"5D",x"66",x"AF",x"66",x"A6",x"66",x"AF",x"AF",x"AF",x"66",x"66",x"A7",x"67",x"66",x"66",x"5E",x"66",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"67",x"67",x"67",x"5F",x"5E",x"5F",x"5F",x"5E",x"5E",x"5E",x"5D",x"15",x"15",x"14",x"5E",x"AF",x"AF",x"AF",x"66",x"5E",x"67",x"66",x"66",x"66",x"65",x"AE",x"65",x"5C",x"5C",x"5C",x"5B",x"53",x"13",x"13",x"0B",x"0B",x"53",x"53",x"53",x"53",x"53",x"53",x"13",x"13",x"13",x"53",x"53",x"5C",x"5C", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"1C",x"1C",x"54",x"53",x"53",x"53",x"53",x"54",x"14",x"1C",x"5C",x"5B",x"5B",x"A3",x"A3",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A2",x"A3",x"9B",x"5C",x"5C",x"65",x"5D",x"66",x"AF",x"AF",x"66",x"66",x"AF",x"6F",x"67",x"66",x"5E",x"67",x"5E",x"67",x"67",x"67",x"AF",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"5E",x"5E",x"67",x"67",x"67",x"67",x"67",x"67",x"5E",x"5D",x"55",x"66",x"AF",x"AF",x"67",x"66",x"5D",x"66",x"66",x"66",x"66",x"5D",x"66",x"65",x"5C",x"5C",x"5C",x"5C",x"5C",x"5C",x"5C",x"5D",x"5C",x"5D",x"5D",x"65",x"65",x"65",x"65",x"65",x"66",x"66",x"AE",x"AE",x"AE",x"AE", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"1C",x"1C",x"5C",x"53",x"53",x"53",x"53",x"53",x"14",x"5C",x"5C",x"5B",x"5B",x"5B",x"A3",x"A3",x"AA",x"A2",x"A2",x"A3",x"A3",x"A3",x"5C",x"5C",x"54",x"5D",x"5D",x"66",x"66",x"66",x"66",x"AF",x"67",x"66",x"5E",x"67",x"5E",x"5E",x"67",x"67",x"66",x"67",x"AF",x"AF",x"AF",x"AF",x"AF",x"A7",x"67",x"67",x"67",x"67",x"5E",x"5E",x"5E",x"5E",x"67",x"67",x"67",x"AF",x"AF",x"67",x"5E",x"5E",x"5E",x"67",x"AF",x"5E",x"A7",x"5E",x"5D",x"5E",x"AF",x"66",x"66",x"66",x"66",x"66",x"66",x"AF",x"AF",x"AF",x"AF",x"AF",x"B7",x"B7",x"B7",x"B7",x"B7",x"B7",x"B7",x"B7",x"B7",x"B7",x"B7",x"B7",x"B7",x"B7",x"B7",x"B7", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"1C",x"1C",x"53",x"53",x"53",x"53",x"53",x"53",x"14",x"54",x"5C",x"5B",x"5B",x"5B",x"A3",x"A3",x"A2",x"A2",x"A2",x"A3",x"A4",x"5C",x"5C",x"5C",x"5D",x"5E",x"5E",x"5D",x"5E",x"66",x"66",x"5E",x"5E",x"5F",x"5E",x"66",x"5E",x"5E",x"67",x"5E",x"67",x"67",x"67",x"A7",x"AF",x"AF",x"AF",x"67",x"67",x"67",x"67",x"67",x"67",x"5E",x"66",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"5E",x"5E",x"AF",x"AF",x"67",x"67",x"5E",x"5E",x"5E",x"66",x"66",x"66",x"66",x"66",x"66",x"66",x"AF",x"B7",x"B7",x"B7",x"B7",x"B7",x"B7",x"B7",x"B7",x"B7",x"AF",x"AF",x"AF",x"AF",x"AF",x"AF",x"AF",x"AF",x"AF",x"AF",x"AF", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"1C",x"14",x"13",x"53",x"53",x"53",x"53",x"53",x"54",x"5C",x"5C",x"5C",x"5B",x"5B",x"A3",x"A3",x"A2",x"A3",x"A3",x"A3",x"A4",x"5B",x"53",x"54",x"5D",x"5D",x"66",x"67",x"67",x"66",x"66",x"5E",x"5E",x"15",x"5E",x"5E",x"67",x"67",x"66",x"67",x"67",x"67",x"67",x"67",x"AF",x"AF",x"A7",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"5E",x"5E",x"67",x"AF",x"67",x"5E",x"67",x"66",x"66",x"5E",x"66",x"AF",x"66",x"66",x"66",x"66",x"AF",x"AF",x"AF",x"AF",x"B7",x"6F",x"6F",x"6F",x"6F",x"B7",x"B7",x"B7",x"B7",x"B7",x"B7",x"B7",x"B7",x"B7",x"B7",x"B7",x"B7", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"14",x"14",x"13",x"53",x"53",x"53",x"53",x"13",x"14",x"14",x"5C",x"5C",x"5B",x"5B",x"A3",x"A3",x"A3",x"A3",x"A3",x"A3",x"A4",x"5B",x"53",x"54",x"5D",x"5D",x"67",x"AF",x"66",x"5D",x"5D",x"5E",x"5E",x"5E",x"5E",x"67",x"B7",x"67",x"67",x"67",x"AF",x"67",x"67",x"67",x"67",x"67",x"67",x"66",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"5E",x"5D",x"5D",x"66",x"6F",x"67",x"5E",x"67",x"67",x"66",x"66",x"6F",x"AF",x"AF",x"AF",x"67",x"66",x"66",x"AF",x"B7",x"B7",x"B7",x"B7",x"77",x"77",x"B7",x"6F",x"6F",x"AF",x"AF",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"1C",x"14",x"53",x"53",x"53",x"53",x"53",x"53",x"13",x"14",x"1C",x"5C",x"5C",x"5C",x"A3",x"A4",x"A3",x"A3",x"A3",x"A3",x"5C",x"53",x"53",x"5C",x"5D",x"66",x"AF",x"66",x"5E",x"66",x"67",x"5E",x"15",x"5E",x"AF",x"67",x"67",x"67",x"66",x"67",x"AF",x"AF",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"66",x"5E",x"66",x"66",x"AF",x"66",x"66",x"5E",x"67",x"5E",x"67",x"AF",x"AF",x"AF",x"AF",x"AF",x"66",x"66",x"67",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"1C",x"14",x"53",x"53",x"53",x"53",x"53",x"53",x"14",x"14",x"14",x"5C",x"5C",x"5B",x"5B",x"63",x"A3",x"A3",x"5C",x"5B",x"5B",x"53",x"54",x"5D",x"66",x"66",x"5E",x"5E",x"67",x"AF",x"67",x"5E",x"16",x"5F",x"67",x"67",x"67",x"5E",x"67",x"67",x"AF",x"AF",x"AF",x"AF",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"6F",x"6F",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"AF",x"67",x"67",x"AF",x"67",x"67",x"5E",x"67",x"5D",x"AF",x"AF",x"AF",x"AF",x"AF",x"AF",x"AF",x"66",x"67",x"AF",x"B7",x"AF",x"6F",x"77",x"B7",x"77",x"B7",x"B7",x"AF",x"B7",x"B7",x"B7",x"B7",x"B7",x"B7",x"B7",x"B7",x"B7", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"14",x"54",x"53",x"53",x"53",x"53",x"53",x"53",x"14",x"14",x"14",x"14",x"5B",x"53",x"5B",x"5B",x"5B",x"5C",x"5C",x"5C",x"5B",x"13",x"54",x"5D",x"66",x"5D",x"5D",x"5E",x"67",x"5E",x"1D",x"1E",x"67",x"56",x"5F",x"5E",x"5E",x"67",x"67",x"AF",x"6F",x"6F",x"6F",x"6F",x"67",x"67",x"67",x"67",x"67",x"67",x"6F",x"67",x"67",x"AF",x"AF",x"6F",x"6F",x"6F",x"6F",x"67",x"67",x"6F",x"AF",x"AF",x"67",x"AF",x"AF",x"A7",x"A7",x"5E",x"67",x"5E",x"67",x"AF",x"67",x"6F",x"AF",x"AF",x"AF",x"67",x"66",x"AF",x"AF",x"AF",x"6F",x"6F",x"77",x"6F",x"B7",x"AF",x"6F",x"6F",x"6F",x"77",x"77",x"77",x"6F",x"AF",x"AF",x"AF", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"54",x"54",x"53",x"53",x"53",x"53",x"53",x"13",x"14",x"14",x"13",x"14",x"5B",x"5B",x"5B",x"5B",x"5C",x"5C",x"5C",x"5C",x"5C",x"13",x"54",x"5D",x"5D",x"5E",x"66",x"5E",x"5E",x"1D",x"5E",x"67",x"5F",x"5E",x"5E",x"56",x"0D",x"67",x"AF",x"67",x"6F",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"AF",x"AF",x"6F",x"6F",x"AF",x"AF",x"AF",x"AF",x"AF",x"67",x"67",x"6F",x"AF",x"AF",x"66",x"66",x"AF",x"67",x"AF",x"67",x"5E",x"67",x"5E",x"67",x"AF",x"66",x"AF",x"AF",x"66",x"AF",x"67",x"66",x"AF",x"B7",x"B7",x"AF",x"77",x"77",x"6F",x"B7",x"6F",x"6F",x"6E",x"6F",x"6F",x"77",x"77",x"77",x"AF",x"AF",x"AF", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"54",x"53",x"53",x"53",x"53",x"53",x"53",x"13",x"13",x"13",x"14",x"14",x"53",x"53",x"5B",x"5C",x"5C",x"5C",x"5C",x"5C",x"13",x"54",x"5D",x"66",x"5D",x"5E",x"5E",x"5E",x"5E",x"66",x"67",x"5E",x"67",x"5F",x"15",x"0D",x"15",x"5F",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"6F",x"AF",x"AF",x"AF",x"AF",x"AF",x"AF",x"AF",x"67",x"67",x"AF",x"AF",x"67",x"67",x"67",x"66",x"AF",x"67",x"AF",x"AF",x"5E",x"5E",x"5E",x"67",x"67",x"67",x"66",x"67",x"AF",x"AF",x"67",x"66",x"6F",x"B7",x"AF",x"AF",x"B7",x"6F",x"B7",x"B7",x"6F",x"6F",x"6E",x"6F",x"B7",x"6F",x"6F",x"77",x"6F",x"AF",x"6F", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"54",x"53",x"53",x"53",x"53",x"53",x"53",x"13",x"13",x"13",x"13",x"54",x"53",x"53",x"5B",x"5C",x"64",x"64",x"5C",x"5C",x"13",x"54",x"5D",x"5E",x"5D",x"67",x"5E",x"15",x"5E",x"67",x"66",x"5E",x"67",x"5E",x"15",x"0C",x"0D",x"56",x"5F",x"67",x"67",x"66",x"66",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"6F",x"AF",x"AF",x"AF",x"AF",x"AF",x"6F",x"67",x"67",x"6F",x"AF",x"67",x"67",x"67",x"66",x"AF",x"67",x"67",x"A7",x"56",x"5E",x"67",x"67",x"66",x"66",x"66",x"67",x"AF",x"A7",x"67",x"66",x"6F",x"B7",x"B7",x"6F",x"B7",x"6F",x"B7",x"6F",x"B7",x"B7",x"6F",x"6F",x"B7",x"6F",x"B7",x"77",x"6F",x"6F",x"6F", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"53",x"53",x"53",x"53",x"53",x"53",x"13",x"13",x"13",x"13",x"13",x"53",x"53",x"53",x"53",x"5C",x"65",x"5C",x"5C",x"53",x"13",x"54",x"55",x"5D",x"5E",x"67",x"5E",x"5D",x"5E",x"66",x"5D",x"66",x"66",x"5E",x"0D",x"0C",x"0D",x"0D",x"56",x"5F",x"5E",x"5E",x"5E",x"5E",x"5E",x"5F",x"5F",x"67",x"67",x"67",x"67",x"67",x"6F",x"AF",x"AF",x"AF",x"67",x"67",x"67",x"6F",x"6F",x"67",x"67",x"67",x"66",x"67",x"67",x"67",x"67",x"56",x"5E",x"67",x"5E",x"5E",x"66",x"66",x"67",x"67",x"67",x"66",x"66",x"66",x"B7",x"B7",x"6F",x"B7",x"6F",x"77",x"6F",x"AF",x"B7",x"6F",x"6F",x"77",x"6F",x"77",x"6F",x"6F",x"6F",x"6F", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"53",x"53",x"53",x"53",x"53",x"13",x"13",x"13",x"13",x"13",x"53",x"53",x"53",x"53",x"53",x"5B",x"64",x"5C",x"5C",x"13",x"54",x"54",x"55",x"5D",x"5E",x"66",x"5E",x"5E",x"5E",x"5D",x"54",x"66",x"5E",x"55",x"0D",x"0D",x"0D",x"0D",x"56",x"5F",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5F",x"5F",x"67",x"67",x"67",x"67",x"6F",x"6F",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"5E",x"67",x"67",x"67",x"67",x"16",x"5E",x"5F",x"5E",x"67",x"67",x"67",x"67",x"67",x"67",x"66",x"66",x"66",x"AF",x"B7",x"6F",x"B7",x"77",x"6F",x"B7",x"6F",x"AF",x"6F",x"6F",x"77",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"53",x"53",x"53",x"53",x"13",x"13",x"13",x"13",x"13",x"13",x"53",x"53",x"53",x"53",x"13",x"5B",x"5C",x"5B",x"5C",x"12",x"54",x"5C",x"5D",x"5D",x"5D",x"5E",x"5E",x"5D",x"5D",x"66",x"5D",x"14",x"5E",x"55",x"0C",x"0D",x"0D",x"0D",x"0D",x"56",x"5F",x"5F",x"67",x"5E",x"5E",x"5E",x"5F",x"5F",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5F",x"5E",x"16",x"56",x"5F",x"5E",x"67",x"67",x"67",x"66",x"66",x"67",x"67",x"66",x"66",x"6F",x"AF",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"67",x"6F",x"6F",x"67",x"6F",x"6F",x"6F",x"6F",x"6F", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"53",x"53",x"13",x"13",x"13",x"13",x"13",x"13",x"53",x"53",x"53",x"53",x"53",x"53",x"53",x"5B",x"5C",x"A4",x"5B",x"53",x"54",x"5C",x"5D",x"5D",x"1D",x"5E",x"5E",x"5D",x"5D",x"5D",x"5C",x"0B",x"5D",x"54",x"0C",x"0D",x"0D",x"0D",x"0D",x"0E",x"5F",x"5F",x"67",x"67",x"67",x"67",x"67",x"5F",x"5F",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"66",x"67",x"67",x"56",x"16",x"16",x"56",x"5E",x"67",x"67",x"67",x"5E",x"66",x"67",x"67",x"66",x"66",x"67",x"67",x"6F",x"6F",x"66",x"66",x"66",x"67",x"67",x"67",x"5E",x"67",x"67",x"6F",x"6F",x"6F",x"6F",x"6F", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"53",x"53",x"13",x"13",x"13",x"13",x"13",x"13",x"53",x"53",x"53",x"53",x"53",x"53",x"53",x"5B",x"5B",x"A4",x"5B",x"53",x"54",x"5C",x"5D",x"1D",x"1D",x"15",x"5E",x"5D",x"5D",x"14",x"13",x"53",x"54",x"54",x"0C",x"0D",x"0D",x"0D",x"0E",x"0E",x"56",x"5E",x"5F",x"67",x"67",x"67",x"67",x"67",x"67",x"5F",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"67",x"67",x"67",x"16",x"16",x"0D",x"0D",x"56",x"5F",x"67",x"5E",x"5E",x"66",x"67",x"67",x"66",x"66",x"5E",x"5E",x"67",x"67",x"1E",x"1E",x"1E",x"5F",x"67",x"5E",x"1E",x"1E",x"1E",x"67",x"6F",x"6F",x"6F",x"6F", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"53",x"53",x"13",x"13",x"13",x"13",x"13",x"13",x"53",x"53",x"53",x"53",x"53",x"53",x"54",x"5B",x"5B",x"AD",x"53",x"53",x"54",x"5C",x"5D",x"1D",x"1D",x"5E",x"5D",x"14",x"66",x"54",x"13",x"0B",x"54",x"54",x"0C",x"0D",x"0D",x"0E",x"0E",x"0E",x"0D",x"56",x"5E",x"5F",x"67",x"67",x"67",x"67",x"67",x"67",x"5F",x"67",x"67",x"67",x"67",x"67",x"67",x"5F",x"5E",x"56",x"16",x"5E",x"5F",x"67",x"67",x"67",x"67",x"5E",x"0D",x"0D",x"16",x"56",x"56",x"5F",x"5F",x"5E",x"5E",x"66",x"67",x"66",x"67",x"67",x"5E",x"5E",x"6F",x"6F",x"1E",x"5F",x"1E",x"5F",x"67",x"5F",x"1F",x"1F",x"1F",x"67",x"6F",x"6F",x"6F",x"6F", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"53",x"53",x"53",x"53",x"13",x"53",x"53",x"53",x"53",x"13",x"13",x"53",x"53",x"53",x"53",x"53",x"53",x"A4",x"53",x"53",x"54",x"55",x"5D",x"5D",x"5E",x"5D",x"15",x"55",x"5D",x"5C",x"13",x"0B",x"54",x"0C",x"0C",x"0C",x"0D",x"0D",x"0E",x"0E",x"0D",x"0D",x"16",x"56",x"5F",x"A7",x"A7",x"A7",x"67",x"67",x"67",x"5F",x"67",x"67",x"67",x"5F",x"67",x"5E",x"56",x"5E",x"5E",x"5E",x"67",x"67",x"A7",x"5F",x"56",x"0D",x"0D",x"0D",x"56",x"57",x"56",x"56",x"56",x"5E",x"5E",x"66",x"66",x"66",x"66",x"67",x"66",x"66",x"67",x"67",x"1E",x"67",x"5F",x"5F",x"67",x"1E",x"67",x"67",x"1E",x"67",x"6F",x"6F",x"6F",x"6F", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"53",x"53",x"53",x"53",x"53",x"53",x"53",x"53",x"53",x"53",x"13",x"53",x"53",x"53",x"53",x"53",x"53",x"64",x"13",x"13",x"54",x"5D",x"5D",x"5D",x"5E",x"5D",x"55",x"55",x"54",x"54",x"54",x"0B",x"0C",x"0C",x"0C",x"0C",x"0D",x"0D",x"0D",x"0E",x"0D",x"0D",x"0D",x"0D",x"56",x"5F",x"A7",x"A7",x"A7",x"67",x"67",x"5F",x"67",x"67",x"67",x"5F",x"5F",x"5E",x"56",x"5E",x"5F",x"5F",x"67",x"67",x"56",x"56",x"0D",x"0D",x"0D",x"0D",x"4E",x"56",x"4E",x"56",x"56",x"5E",x"5E",x"66",x"66",x"66",x"66",x"67",x"5E",x"66",x"67",x"67",x"1E",x"5F",x"5F",x"5F",x"67",x"1E",x"67",x"67",x"1E",x"67",x"6F",x"6F",x"6F",x"6F", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"53",x"53",x"53",x"53",x"53",x"53",x"53",x"53",x"53",x"53",x"53",x"53",x"53",x"53",x"53",x"53",x"53",x"5C",x"13",x"13",x"54",x"55",x"5D",x"5D",x"5E",x"55",x"5D",x"14",x"0B",x"54",x"54",x"0B",x"0C",x"0C",x"0C",x"0D",x"0D",x"0D",x"0E",x"0E",x"0E",x"0E",x"0E",x"0D",x"0D",x"0D",x"16",x"56",x"5F",x"5F",x"5F",x"5F",x"5F",x"67",x"5F",x"5F",x"5E",x"56",x"15",x"15",x"16",x"16",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0E",x"0E",x"0E",x"0E",x"0E",x"56",x"56",x"5E",x"5E",x"67",x"66",x"66",x"67",x"67",x"5E",x"5E",x"67",x"67",x"1E",x"1E",x"1E",x"5F",x"67",x"1E",x"27",x"67",x"5E",x"67",x"6F",x"6F",x"6F",x"6F", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"53",x"53",x"53",x"53",x"53",x"53",x"53",x"53",x"53",x"53",x"53",x"53",x"53",x"53",x"53",x"53",x"13",x"53",x"13",x"13",x"54",x"55",x"5D",x"5D",x"5E",x"5D",x"55",x"14",x"0B",x"54",x"54",x"0B",x"0C",x"0C",x"0C",x"0D",x"0D",x"0D",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0E",x"0D",x"0D",x"0D",x"0E",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"16",x"56",x"5E",x"5F",x"67",x"66",x"66",x"67",x"67",x"5E",x"1E",x"26",x"67",x"1E",x"1E",x"1E",x"5E",x"67",x"1E",x"27",x"67",x"1E",x"67",x"6F",x"6F",x"6F",x"6F", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"13",x"13",x"53",x"53",x"53",x"53",x"53",x"53",x"53",x"53",x"53",x"53",x"53",x"53",x"53",x"53",x"53",x"53",x"13",x"13",x"54",x"55",x"5D",x"5E",x"5D",x"5D",x"15",x"14",x"54",x"54",x"13",x"0B",x"0C",x"0C",x"0C",x"0D",x"0D",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0D",x"0D",x"0D",x"0D",x"0E",x"0E",x"0E",x"0E",x"4E",x"0E",x"0D",x"0D",x"0E",x"0E",x"0E",x"0E",x"4E",x"0E",x"56",x"56",x"5E",x"5E",x"66",x"66",x"66",x"67",x"67",x"5E",x"1E",x"1E",x"67",x"1E",x"5F",x"5E",x"1E",x"67",x"1E",x"1E",x"1E",x"1E",x"67",x"67",x"6F",x"6F",x"6F", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"13",x"13",x"53",x"53",x"53",x"53",x"53",x"53",x"53",x"53",x"53",x"53",x"13",x"13",x"53",x"53",x"53",x"13",x"13",x"13",x"54",x"55",x"5D",x"5E",x"55",x"5D",x"15",x"14",x"54",x"53",x"0B",x"53",x"0C",x"0C",x"0C",x"01",x"0D",x"0D",x"0E",x"0E",x"4E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"4E",x"4E",x"4E",x"0E",x"0E",x"0D",x"0D",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"56",x"5E",x"5E",x"66",x"66",x"67",x"67",x"67",x"66",x"66",x"1E",x"27",x"1E",x"67",x"67",x"1E",x"67",x"1E",x"1E",x"1D",x"5E",x"67",x"6F",x"6F",x"6F",x"6F", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"13",x"13",x"53",x"53",x"53",x"53",x"53",x"53",x"53",x"53",x"53",x"13",x"13",x"13",x"53",x"53",x"53",x"0B",x"53",x"14",x"5D",x"55",x"5D",x"5D",x"55",x"5D",x"55",x"54",x"54",x"0B",x"0B",x"53",x"0C",x"0C",x"0C",x"01",x"0D",x"0D",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"4E",x"0E",x"0E",x"0E",x"4E",x"4E",x"0E",x"4E",x"4E",x"4E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"56",x"56",x"5E",x"5E",x"67",x"67",x"67",x"67",x"67",x"67",x"27",x"67",x"67",x"67",x"67",x"67",x"67",x"26",x"26",x"1E",x"66",x"67",x"6F",x"6F",x"6F",x"6F", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"13",x"13",x"53",x"53",x"53",x"53",x"53",x"53",x"53",x"53",x"53",x"53",x"13",x"53",x"53",x"53",x"53",x"0B",x"54",x"54",x"5D",x"55",x"5D",x"15",x"5D",x"55",x"5D",x"55",x"0B",x"0B",x"13",x"0B",x"0C",x"0C",x"0C",x"0C",x"0D",x"0D",x"0D",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"4E",x"0E",x"0D",x"0D",x"16",x"56",x"5E",x"5E",x"67",x"67",x"67",x"67",x"67",x"6F",x"6F",x"6F",x"67",x"6F",x"67",x"67",x"6F",x"67",x"6F",x"6F",x"6F",x"67",x"66",x"66",x"AE",x"B7", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"13",x"13",x"13",x"53",x"53",x"53",x"53",x"53",x"53",x"53",x"53",x"53",x"13",x"13",x"13",x"53",x"53",x"13",x"13",x"54",x"5D",x"5D",x"5D",x"15",x"5D",x"5D",x"5D",x"14",x"0B",x"0B",x"13",x"0B",x"0B",x"0C",x"0C",x"0C",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0D",x"15",x"56",x"5E",x"66",x"67",x"67",x"67",x"67",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"5E",x"14",x"53",x"5B",x"A5",x"07", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"13",x"13",x"13",x"53",x"53",x"53",x"53",x"53",x"53",x"53",x"53",x"53",x"13",x"53",x"53",x"53",x"53",x"13",x"13",x"54",x"5D",x"5D",x"5D",x"15",x"5D",x"5D",x"5D",x"14",x"0B",x"0B",x"4B",x"0B",x"0B",x"0C",x"0C",x"0C",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0D",x"0D",x"15",x"56",x"5E",x"66",x"66",x"67",x"67",x"67",x"67",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"67",x"6F",x"6F",x"6F",x"66",x"5D",x"5C",x"5B",x"5B",x"5C", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"53",x"13",x"13",x"53",x"53",x"53",x"53",x"53",x"53",x"53",x"53",x"53",x"13",x"13",x"13",x"53",x"53",x"13",x"13",x"54",x"5D",x"5D",x"5D",x"55",x"55",x"5D",x"5D",x"14",x"0B",x"0B",x"0B",x"0B",x"0B",x"0C",x"0C",x"0C",x"0C",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"15",x"56",x"5E",x"66",x"66",x"67",x"67",x"67",x"67",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"67",x"67",x"6F",x"6F",x"67",x"66",x"5C",x"14",x"14",x"5C", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"13",x"13",x"13",x"53",x"53",x"53",x"53",x"53",x"53",x"53",x"53",x"53",x"13",x"13",x"13",x"13",x"53",x"13",x"13",x"54",x"5D",x"5D",x"5D",x"5D",x"55",x"5D",x"5D",x"14",x"0B",x"0B",x"0B",x"0B",x"0B",x"0C",x"0C",x"0C",x"0C",x"0C",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"15",x"56",x"5E",x"5E",x"67",x"67",x"67",x"66",x"67",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"67",x"6F",x"6F",x"6F",x"67",x"66",x"66",x"66",x"66", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"13",x"13",x"13",x"53",x"53",x"53",x"53",x"53",x"53",x"53",x"53",x"53",x"13",x"13",x"13",x"13",x"53",x"13",x"13",x"54",x"5D",x"5D",x"5D",x"5E",x"5D",x"5E",x"5D",x"55",x"0B",x"0B",x"0B",x"0B",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"01",x"0C",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"15",x"55",x"5E",x"5E",x"67",x"67",x"67",x"66",x"67",x"6F",x"6F",x"6F",x"6F",x"67",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"67",x"6F",x"6F",x"67",x"67", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"13",x"13",x"13",x"13",x"53",x"53",x"53",x"52",x"52",x"52",x"53",x"53",x"53",x"13",x"13",x"13",x"13",x"13",x"13",x"54",x"5D",x"5D",x"5D",x"5E",x"5E",x"5E",x"5E",x"55",x"0B",x"0B",x"0B",x"0B",x"0C",x"0C",x"0C",x"0C",x"01",x"01",x"01",x"01",x"0C",x"0C",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"15",x"55",x"5E",x"5E",x"67",x"67",x"66",x"66",x"67",x"6F",x"6F",x"6F",x"6F",x"67",x"67",x"6F",x"6F",x"6F",x"6F",x"67",x"67",x"67",x"67",x"67",x"67",x"67", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"13",x"13",x"13",x"13",x"53",x"53",x"52",x"12",x"12",x"12",x"53",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"54",x"5D",x"5D",x"5D",x"5E",x"5E",x"5E",x"5E",x"55",x"0C",x"0B",x"0B",x"0B",x"0C",x"0C",x"0C",x"0C",x"01",x"01",x"01",x"01",x"0C",x"0C",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"15",x"15",x"55",x"5E",x"66",x"67",x"66",x"66",x"67",x"6F",x"6F",x"6F",x"6F",x"67",x"67",x"67",x"6F",x"6F",x"6F",x"67",x"67",x"67",x"67",x"67",x"6F",x"6F", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"13",x"13",x"13",x"13",x"53",x"53",x"52",x"12",x"12",x"12",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"54",x"5D",x"5D",x"5E",x"5E",x"5E",x"5E",x"5E",x"55",x"0C",x"0B",x"0B",x"0B",x"0C",x"0C",x"0C",x"0C",x"01",x"01",x"01",x"01",x"0C",x"0C",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"15",x"15",x"55",x"5E",x"66",x"67",x"66",x"66",x"67",x"6F",x"6F",x"6F",x"6F",x"67",x"67",x"67",x"67",x"6F",x"6F",x"67",x"67",x"67",x"6F",x"6F",x"67",x"67", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"13",x"13",x"13",x"13",x"53",x"53",x"52",x"52",x"52",x"52",x"12",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"14",x"55",x"5D",x"5E",x"5E",x"5E",x"5F",x"5E",x"5E",x"54",x"0B",x"0B",x"0B",x"0C",x"0C",x"0C",x"0C",x"01",x"01",x"0C",x"0D",x"0C",x"0C",x"0C",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"01",x"0D",x"0D",x"0D",x"4D",x"0C",x"54",x"0C",x"54",x"15",x"5E",x"66",x"67",x"67",x"66",x"66",x"67",x"6F",x"67",x"67",x"67",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"67",x"67",x"67",x"67",x"67",x"67", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"13",x"13",x"13",x"13",x"53",x"53",x"52",x"52",x"12",x"12",x"12",x"12",x"53",x"13",x"13",x"13",x"53",x"13",x"13",x"54",x"55",x"5E",x"5E",x"5E",x"5E",x"5F",x"5F",x"5E",x"55",x"54",x"0B",x"0B",x"0C",x"0C",x"0C",x"0C",x"01",x"01",x"0C",x"0D",x"0C",x"0C",x"0C",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"01",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"4D",x"0C",x"0B",x"0B",x"14",x"15",x"5E",x"5E",x"67",x"67",x"66",x"66",x"67",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"67",x"67",x"67",x"67", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"13",x"13",x"13",x"13",x"13",x"12",x"52",x"52",x"12",x"12",x"12",x"53",x"53",x"53",x"13",x"13",x"53",x"13",x"13",x"54",x"55",x"5E",x"5E",x"5E",x"5E",x"67",x"5F",x"5E",x"5D",x"5D",x"0B",x"0C",x"0C",x"0C",x"0C",x"0C",x"01",x"01",x"0D",x"0D",x"0C",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"56",x"55",x"0B",x"0B",x"0C",x"15",x"5E",x"5E",x"66",x"67",x"66",x"66",x"6F",x"AF",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"13",x"13",x"13",x"13",x"13",x"12",x"52",x"52",x"12",x"12",x"12",x"53",x"53",x"53",x"13",x"13",x"53",x"13",x"13",x"14",x"55",x"5E",x"5E",x"5E",x"5E",x"67",x"5F",x"5E",x"5D",x"5D",x"0B",x"0C",x"0C",x"0C",x"0C",x"0C",x"01",x"01",x"01",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0E",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"56",x"66",x"0B",x"14",x"0B",x"15",x"5E",x"5E",x"66",x"A6",x"66",x"66",x"6F",x"AF",x"B7",x"77",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"13",x"13",x"13",x"12",x"12",x"12",x"52",x"52",x"12",x"12",x"12",x"53",x"53",x"53",x"13",x"13",x"13",x"0B",x"13",x"14",x"55",x"5E",x"5E",x"5E",x"5E",x"67",x"67",x"5E",x"54",x"5D",x"0B",x"0C",x"0C",x"0C",x"0C",x"01",x"01",x"01",x"01",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0E",x"0E",x"0E",x"56",x"AF",x"13",x"14",x"0B",x"14",x"5E",x"5E",x"66",x"66",x"66",x"66",x"66",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"13",x"13",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"12",x"53",x"53",x"53",x"53",x"13",x"13",x"0B",x"13",x"13",x"55",x"5E",x"5E",x"5E",x"67",x"67",x"67",x"5E",x"54",x"5C",x"0B",x"0B",x"0C",x"0C",x"0C",x"01",x"01",x"01",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"56",x"AF",x"14",x"0B",x"0B",x"14",x"5D",x"5E",x"66",x"66",x"66",x"66",x"66",x"67",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"13",x"13",x"12",x"12",x"12",x"12",x"52",x"52",x"52",x"12",x"12",x"52",x"53",x"53",x"53",x"13",x"13",x"0B",x"13",x"13",x"55",x"5E",x"5E",x"5E",x"67",x"67",x"67",x"5E",x"54",x"5C",x"54",x"0B",x"0C",x"0C",x"0C",x"01",x"01",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"5E",x"AF",x"5D",x"0B",x"0B",x"14",x"5D",x"5E",x"66",x"67",x"67",x"67",x"67",x"67",x"67",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"13",x"13",x"12",x"12",x"12",x"12",x"52",x"52",x"52",x"52",x"12",x"12",x"53",x"53",x"53",x"13",x"13",x"0B",x"13",x"13",x"55",x"5E",x"5E",x"5E",x"67",x"5F",x"67",x"66",x"5C",x"5C",x"5C",x"0B",x"0C",x"0C",x"0C",x"0C",x"01",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"56",x"56",x"16",x"0E",x"0E",x"5E",x"AF",x"66",x"0B",x"0B",x"0C",x"55",x"5E",x"66",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F",x"6F", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"13",x"13",x"12",x"12",x"12",x"12",x"52",x"52",x"12",x"52",x"52",x"52",x"53",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"55",x"5E",x"5E",x"67",x"67",x"5E",x"5F",x"5E",x"5C",x"54",x"54",x"54",x"0C",x"0C",x"0C",x"01",x"01",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0E",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"56",x"57",x"5F",x"56",x"56",x"57",x"5F",x"57",x"5E",x"AF",x"66",x"14",x"0B",x"0C",x"15",x"5E",x"5E",x"5F",x"5E",x"67",x"67",x"5E",x"67",x"6F",x"67",x"6F",x"6F",x"67",x"6F",x"6F",x"6F",x"6F",x"6F",x"67",x"6F",x"6F",x"6F", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"13",x"13",x"12",x"12",x"12",x"12",x"52",x"52",x"12",x"52",x"52",x"52",x"53",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"55",x"5E",x"5E",x"67",x"67",x"66",x"5F",x"5E",x"5C",x"5C",x"5C",x"54",x"0B",x"0C",x"0C",x"01",x"01",x"01",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"01",x"0E",x"0D",x"0D",x"0D",x"56",x"56",x"57",x"0E",x"0D",x"0D",x"0D",x"0D",x"0E",x"67",x"5E",x"5E",x"5D",x"13",x"0B",x"14",x"55",x"5E",x"66",x"5E",x"5E",x"67",x"67",x"67",x"66",x"66",x"66",x"66",x"66",x"66",x"66",x"66",x"66",x"67",x"6F",x"67",x"67",x"6F",x"6F", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"13",x"13",x"12",x"12",x"12",x"52",x"52",x"52",x"52",x"52",x"52",x"52",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"55",x"5E",x"5E",x"67",x"67",x"67",x"5E",x"5E",x"5C",x"5C",x"5C",x"5C",x"0C",x"0C",x"0C",x"0C",x"0D",x"01",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0E",x"0D",x"0D",x"0D",x"57",x"16",x"0D",x"0D",x"56",x"56",x"5E",x"5F",x"56",x"5F",x"16",x"0C",x"13",x"0B",x"0C",x"55",x"5D",x"5E",x"66",x"66",x"66",x"66",x"66",x"66",x"5D",x"14",x"14",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"14",x"14",x"14",x"14", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"12",x"12",x"12",x"12",x"52",x"52",x"52",x"52",x"52",x"52",x"52",x"52",x"52",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"5D",x"5E",x"67",x"67",x"67",x"66",x"5E",x"5E",x"5C",x"5B",x"5C",x"54",x"54",x"0C",x"0C",x"0C",x"0D",x"01",x"01",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0E",x"0D",x"0D",x"0D",x"56",x"56",x"56",x"16",x"5E",x"67",x"AF",x"5E",x"5E",x"16",x"0D",x"67",x"0B",x"0B",x"0B",x"0B",x"55",x"5D",x"5E",x"66",x"66",x"66",x"66",x"66",x"A6",x"5D",x"13",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"12",x"12",x"0A",x"0A",x"0A",x"0A", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"12",x"12",x"12",x"12",x"52",x"52",x"52",x"52",x"52",x"52",x"12",x"52",x"12",x"12",x"13",x"13",x"13",x"13",x"13",x"13",x"5D",x"5E",x"67",x"67",x"67",x"66",x"5E",x"5D",x"5C",x"53",x"53",x"53",x"54",x"0C",x"0B",x"0C",x"0D",x"0D",x"01",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"5F",x"5F",x"67",x"67",x"A7",x"5E",x"5E",x"5E",x"0D",x"16",x"15",x"5E",x"14",x"0B",x"0B",x"0B",x"55",x"5E",x"66",x"66",x"A7",x"5E",x"66",x"A6",x"A6",x"A6",x"5D",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"0A",x"0A",x"0A",x"12",x"12",x"52",x"52",x"52",x"52",x"52",x"52",x"12",x"12",x"12",x"13",x"13",x"13",x"13",x"13",x"13",x"5D",x"5F",x"67",x"67",x"67",x"66",x"5E",x"5D",x"5C",x"53",x"53",x"53",x"54",x"0B",x"0B",x"0C",x"0C",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"5F",x"5F",x"5F",x"5E",x"15",x"5E",x"6F",x"AF",x"5E",x"0D",x"0D",x"5F",x"55",x"54",x"54",x"0B",x"55",x"5E",x"66",x"67",x"67",x"5E",x"66",x"66",x"66",x"AE",x"65",x"12",x"0A",x"0A",x"52",x"52",x"52",x"49",x"51",x"51",x"0A",x"0A",x"0A",x"0A", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"0A",x"0A",x"0A",x"12",x"12",x"52",x"52",x"52",x"52",x"52",x"4A",x"0A",x"0A",x"12",x"13",x"13",x"13",x"13",x"0B",x"13",x"5D",x"5F",x"67",x"67",x"67",x"67",x"5E",x"5D",x"5C",x"5B",x"5B",x"53",x"54",x"0C",x"0B",x"0C",x"0C",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"4E",x"0D",x"0D",x"56",x"5F",x"56",x"15",x"15",x"15",x"67",x"6F",x"AF",x"AF",x"5E",x"0D",x"5F",x"55",x"5D",x"5D",x"0C",x"55",x"5E",x"66",x"67",x"67",x"5F",x"5E",x"66",x"66",x"66",x"65",x"13",x"12",x"52",x"53",x"53",x"52",x"52",x"52",x"52",x"52",x"52",x"52",x"52", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"0A",x"0A",x"0A",x"0A",x"12",x"52",x"52",x"52",x"52",x"52",x"4A",x"0A",x"0A",x"12",x"12",x"13",x"13",x"13",x"0B",x"13",x"5D",x"5F",x"67",x"67",x"67",x"67",x"5E",x"5E",x"5C",x"5B",x"5B",x"5B",x"54",x"54",x"0C",x"0C",x"0C",x"0C",x"0D",x"01",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"5F",x"56",x"0D",x"0D",x"67",x"AF",x"5D",x"AF",x"AF",x"AF",x"A7",x"55",x"5E",x"55",x"5D",x"A6",x"54",x"55",x"5D",x"66",x"67",x"67",x"67",x"5E",x"5E",x"67",x"66",x"65",x"65",x"13",x"53",x"5B",x"5B",x"5B",x"5B",x"5A",x"5A",x"5A",x"52",x"52",x"52", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"52",x"0A",x"0A",x"0A",x"0A",x"0A",x"12",x"52",x"52",x"0A",x"0A",x"12",x"53",x"12",x"12",x"12",x"53",x"0B",x"0B",x"13",x"55",x"5E",x"67",x"67",x"67",x"67",x"5E",x"5E",x"5C",x"5B",x"5B",x"53",x"54",x"54",x"54",x"0B",x"0C",x"0C",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0E",x"0D",x"5F",x"5F",x"0D",x"15",x"5E",x"5E",x"AE",x"AE",x"AF",x"B7",x"AF",x"56",x"5E",x"55",x"55",x"5E",x"5E",x"55",x"5D",x"67",x"66",x"67",x"67",x"66",x"66",x"66",x"66",x"66",x"65",x"53",x"53",x"5B",x"5B",x"52",x"5B",x"5A",x"5A",x"5A",x"5B",x"5B",x"5B", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"52",x"0A",x"0A",x"0A",x"0A",x"0A",x"12",x"12",x"52",x"0A",x"0A",x"12",x"52",x"12",x"12",x"12",x"53",x"0B",x"0B",x"13",x"55",x"5E",x"67",x"67",x"67",x"67",x"5E",x"5E",x"5C",x"5B",x"5C",x"53",x"53",x"54",x"53",x"0B",x"0C",x"0C",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0E",x"0E",x"0D",x"56",x"A7",x"15",x"AF",x"5E",x"5D",x"5D",x"AF",x"AF",x"AF",x"A7",x"15",x"5F",x"15",x"56",x"5E",x"5E",x"55",x"55",x"5E",x"66",x"67",x"66",x"66",x"66",x"66",x"66",x"66",x"65",x"54",x"12",x"12",x"52",x"52",x"52",x"52",x"52",x"52",x"52",x"52",x"52", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"4A",x"0A",x"0A",x"0A",x"0A",x"0A",x"12",x"12",x"52",x"0A",x"0A",x"12",x"52",x"52",x"12",x"12",x"53",x"0B",x"0B",x"13",x"55",x"5E",x"67",x"67",x"67",x"67",x"66",x"5E",x"5C",x"53",x"5B",x"53",x"53",x"53",x"53",x"0B",x"0C",x"0C",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0E",x"0D",x"A7",x"0D",x"55",x"67",x"55",x"0B",x"5D",x"5E",x"5E",x"67",x"5E",x"67",x"15",x"5E",x"67",x"67",x"5E",x"55",x"5E",x"5E",x"66",x"66",x"5E",x"5E",x"66",x"66",x"66",x"65",x"5C",x"0A",x"0A",x"0A",x"52",x"52",x"51",x"52",x"52",x"52",x"52",x"51", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"4A",x"0A",x"0A",x"0A",x"0A",x"0A",x"12",x"12",x"12",x"12",x"0A",x"12",x"12",x"52",x"12",x"12",x"13",x"0B",x"13",x"13",x"55",x"5E",x"67",x"67",x"67",x"67",x"66",x"5D",x"5C",x"53",x"53",x"53",x"53",x"53",x"54",x"0B",x"0B",x"0C",x"0C",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0E",x"0D",x"01",x"5F",x"67",x"0D",x"0D",x"5D",x"AF",x"AF",x"A7",x"AF",x"5E",x"56",x"67",x"15",x"5F",x"67",x"67",x"5E",x"5D",x"5D",x"5E",x"5E",x"5E",x"5E",x"5E",x"66",x"66",x"66",x"66",x"5D",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"52",x"52",x"4A",x"0A",x"0A", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"12",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"12",x"12",x"12",x"0A",x"0A",x"0A",x"12",x"12",x"12",x"13",x"0B",x"13",x"14",x"55",x"5E",x"5F",x"67",x"67",x"67",x"5E",x"5D",x"54",x"53",x"5B",x"53",x"53",x"53",x"54",x"53",x"0B",x"0C",x"0C",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0E",x"0D",x"0E",x"0E",x"0D",x"0D",x"0D",x"5F",x"A7",x"56",x"A7",x"5D",x"55",x"5E",x"0D",x"5E",x"67",x"15",x"5E",x"67",x"67",x"67",x"66",x"5E",x"15",x"5D",x"5E",x"5E",x"5E",x"5E",x"5E",x"66",x"66",x"66",x"5D",x"13",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"12",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"12",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"12",x"0A",x"13",x"0B",x"13",x"54",x"55",x"5E",x"5E",x"67",x"67",x"67",x"5E",x"5D",x"53",x"53",x"53",x"53",x"53",x"53",x"53",x"53",x"0B",x"0C",x"0C",x"0C",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0E",x"0E",x"0E",x"01",x"0E",x"56",x"0D",x"0D",x"5F",x"A7",x"5E",x"56",x"5E",x"56",x"5F",x"A7",x"56",x"15",x"5F",x"67",x"67",x"67",x"67",x"5E",x"15",x"5D",x"5E",x"5E",x"5E",x"5E",x"5E",x"66",x"66",x"66",x"66",x"54",x"14",x"0B",x"0B",x"13",x"53",x"54",x"53",x"14",x"13",x"13", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"0B",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"12",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0B",x"0B",x"13",x"54",x"55",x"5E",x"5E",x"67",x"67",x"67",x"5E",x"55",x"0B",x"12",x"53",x"53",x"53",x"53",x"53",x"53",x"0B",x"0C",x"0C",x"0C",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0E",x"0E",x"0D",x"0D",x"4E",x"01",x"0D",x"4E",x"0D",x"0E",x"5F",x"67",x"A7",x"5F",x"56",x"16",x"0D",x"16",x"67",x"67",x"67",x"67",x"67",x"5E",x"5D",x"1D",x"5E",x"5E",x"5E",x"5E",x"5E",x"66",x"66",x"66",x"66",x"5D",x"5D",x"54",x"13",x"54",x"5C",x"5D",x"66",x"66",x"66",x"66", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"0B",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"12",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0B",x"0B",x"13",x"54",x"5D",x"5E",x"5E",x"67",x"67",x"67",x"66",x"55",x"0A",x"0A",x"0A",x"52",x"52",x"53",x"53",x"53",x"0B",x"0B",x"0C",x"0C",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0E",x"0D",x"0E",x"0D",x"0D",x"4E",x"0D",x"0D",x"0D",x"0D",x"16",x"16",x"0D",x"16",x"56",x"67",x"67",x"67",x"67",x"67",x"66",x"5D",x"5D",x"5D",x"5E",x"5E",x"5E",x"5E",x"66",x"66",x"66",x"66",x"5D",x"5E",x"5D",x"14",x"13",x"13",x"1C",x"5D",x"1E",x"5E",x"5E", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"13",x"13",x"0A",x"0A",x"13",x"13",x"12",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0B",x"0B",x"13",x"54",x"5D",x"5E",x"5E",x"67",x"67",x"67",x"66",x"5D",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"4B",x"0B",x"0B",x"0C",x"0C",x"0C",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0E",x"0D",x"0E",x"0D",x"0D",x"0D",x"0D",x"5F",x"67",x"67",x"67",x"67",x"66",x"66",x"5E",x"5E",x"5D",x"5D",x"5E",x"5E",x"5E",x"5E",x"66",x"66",x"66",x"5E",x"5E",x"5D",x"5D",x"14",x"14",x"14",x"15",x"1E",x"1E",x"1E", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"13",x"13",x"0A",x"0A",x"13",x"13",x"12",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0B",x"0B",x"13",x"54",x"5D",x"5E",x"5E",x"67",x"67",x"67",x"67",x"5D",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0B",x"54",x"0C",x"0C",x"0C",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"4E",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0E",x"0E",x"0E",x"0E",x"0D",x"0D",x"0D",x"15",x"67",x"67",x"67",x"67",x"67",x"66",x"66",x"5E",x"5E",x"5D",x"5D",x"5E",x"5E",x"5E",x"5E",x"66",x"67",x"66",x"5E",x"5E",x"5E",x"5D",x"1D",x"14",x"14",x"14",x"15",x"1D",x"1E", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"13",x"13",x"0B",x"0B",x"13",x"13",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0B",x"0B",x"13",x"54",x"5E",x"5E",x"5E",x"67",x"67",x"67",x"66",x"5D",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0B",x"54",x"55",x"15",x"0C",x"0C",x"0D",x"0D",x"0D",x"0D",x"0D",x"4E",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0E",x"0D",x"0D",x"0E",x"0D",x"0D",x"0D",x"56",x"A7",x"A7",x"A7",x"67",x"67",x"67",x"66",x"5E",x"5E",x"5D",x"5D",x"5D",x"5E",x"5E",x"5E",x"5E",x"67",x"66",x"5E",x"5E",x"5D",x"5D",x"5D",x"1C",x"14",x"13",x"14",x"14",x"1D", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"13",x"13",x"0B",x"0B",x"13",x"13",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0B",x"0B",x"13",x"54",x"5E",x"5E",x"5E",x"67",x"67",x"67",x"66",x"5D",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0B",x"54",x"5D",x"5E",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0E",x"0E",x"0D",x"0D",x"55",x"5E",x"A7",x"A7",x"A7",x"67",x"67",x"67",x"66",x"66",x"5E",x"5E",x"5D",x"1D",x"5D",x"5E",x"5E",x"5E",x"67",x"66",x"5E",x"5D",x"5D",x"5D",x"5D",x"5D",x"5C",x"14",x"13",x"13",x"13", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"13",x"13",x"0B",x"0B",x"0B",x"0B",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0B",x"0B",x"13",x"54",x"5E",x"5E",x"5E",x"67",x"67",x"67",x"66",x"5D",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0B",x"0B",x"55",x"5E",x"5E",x"15",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0E",x"0D",x"0D",x"0D",x"55",x"5E",x"A7",x"A7",x"67",x"67",x"67",x"67",x"67",x"66",x"5E",x"5E",x"5D",x"15",x"5D",x"5D",x"5E",x"5E",x"66",x"66",x"5E",x"5D",x"5D",x"5C",x"5C",x"5C",x"5C",x"5C",x"53",x"13",x"13", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"13",x"13",x"0B",x"0B",x"0B",x"0B",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0B",x"0B",x"13",x"54",x"5E",x"5E",x"5E",x"66",x"67",x"67",x"66",x"55",x"0A",x"0A",x"0A",x"0A",x"4A",x"0A",x"0A",x"0A",x"0B",x"0B",x"14",x"5D",x"5E",x"5E",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0E",x"0D",x"0D",x"0D",x"55",x"67",x"A7",x"A7",x"67",x"67",x"67",x"67",x"67",x"67",x"66",x"66",x"5D",x"55",x"55",x"5D",x"5D",x"5E",x"5E",x"66",x"66",x"5D",x"14",x"13",x"13",x"13",x"13",x"53",x"52",x"52",x"52", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"13",x"13",x"13",x"0B",x"0B",x"0B",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0B",x"0B",x"13",x"54",x"5E",x"5E",x"5E",x"66",x"67",x"67",x"5E",x"54",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0B",x"0B",x"14",x"55",x"5E",x"5E",x"5E",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0E",x"0D",x"0D",x"0D",x"56",x"A7",x"A7",x"67",x"67",x"66",x"67",x"67",x"67",x"67",x"67",x"66",x"5E",x"5D",x"55",x"55",x"5D",x"5E",x"5E",x"5E",x"66",x"5D",x"14",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"13",x"13",x"0B",x"0B",x"0B",x"0B",x"0B",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0B",x"13",x"54",x"5E",x"5E",x"5E",x"5E",x"67",x"66",x"5E",x"54",x"0A",x"0A",x"0A",x"0A",x"00",x"0A",x"0A",x"0A",x"0A",x"0B",x"14",x"55",x"5D",x"5E",x"67",x"56",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0E",x"0D",x"0D",x"0D",x"56",x"A7",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"66",x"5E",x"5D",x"55",x"55",x"5D",x"5E",x"5E",x"5E",x"66",x"5D",x"53",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"13",x"13",x"13",x"13",x"0B",x"0B",x"0B",x"0B",x"0B",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0B",x"13",x"54",x"5E",x"5E",x"5E",x"5E",x"66",x"67",x"66",x"0C",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0B",x"0B",x"13",x"54",x"5D",x"5E",x"5E",x"5F",x"56",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0E",x"0E",x"0D",x"0D",x"0D",x"5F",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"66",x"5E",x"66",x"14",x"14",x"55",x"5E",x"5D",x"66",x"5D",x"5D",x"54",x"0A",x"0A",x"0A",x"00",x"00",x"00",x"00",x"00", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"13",x"13",x"13",x"13",x"0B",x"0B",x"0B",x"0B",x"0B",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0B",x"13",x"54",x"5D",x"5E",x"5E",x"5E",x"66",x"67",x"66",x"0B",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0B",x"0B",x"0B",x"54",x"5D",x"5D",x"5E",x"5F",x"5E",x"16",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0E",x"0E",x"0D",x"0D",x"0D",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"66",x"66",x"66",x"66",x"5D",x"14",x"55",x"5D",x"5D",x"5E",x"5D",x"66",x"5C",x"0A",x"0A",x"0A",x"00",x"00",x"00",x"00",x"00", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"13",x"13",x"13",x"13",x"13",x"0B",x"0B",x"0B",x"0B",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0B",x"0B",x"14",x"5D",x"5E",x"5E",x"66",x"67",x"67",x"5E",x"0B",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0B",x"0B",x"0B",x"14",x"55",x"55",x"5E",x"5E",x"5F",x"5E",x"15",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0E",x"0E",x"0D",x"0D",x"15",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"66",x"66",x"5E",x"5E",x"14",x"14",x"55",x"5D",x"5E",x"5E",x"66",x"5D",x"0A",x"0A",x"0A",x"00",x"00",x"00",x"00",x"00", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"0B",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0B",x"13",x"55",x"5E",x"5E",x"67",x"67",x"67",x"5E",x"0B",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0B",x"0B",x"0B",x"14",x"55",x"5D",x"5D",x"5E",x"5E",x"5F",x"5E",x"15",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0E",x"0D",x"0D",x"0D",x"55",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"67",x"66",x"A7",x"5E",x"66",x"55",x"14",x"15",x"5D",x"5D",x"5E",x"66",x"5D",x"0B",x"0A",x"00",x"00",x"00",x"00",x"00",x"00", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"13",x"13",x"13",x"13",x"12",x"12",x"12",x"12",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"13",x"55",x"5E",x"5E",x"67",x"67",x"67",x"5E",x"0B",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0B",x"0B",x"0B",x"0B",x"54",x"55",x"5D",x"5E",x"5E",x"5E",x"5E",x"5E",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0E",x"0D",x"0D",x"0D",x"56",x"67",x"67",x"67",x"66",x"66",x"66",x"67",x"67",x"67",x"67",x"67",x"A7",x"A7",x"66",x"66",x"5D",x"0C",x"15",x"55",x"5D",x"5E",x"66",x"5D",x"53",x"0A",x"0A",x"00",x"00",x"00",x"00",x"00", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"13",x"13",x"13",x"13",x"12",x"12",x"12",x"12",x"12",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"13",x"55",x"5E",x"5E",x"66",x"66",x"66",x"5E",x"0B",x"0A",x"0A",x"00",x"0A",x"0A",x"0A",x"0A",x"0A",x"0B",x"0B",x"0B",x"0B",x"14",x"55",x"5D",x"5E",x"5E",x"5E",x"5E",x"5F",x"56",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"5E",x"67",x"67",x"66",x"66",x"66",x"66",x"66",x"67",x"67",x"67",x"67",x"A7",x"66",x"66",x"5E",x"5E",x"14",x"14",x"15",x"5D",x"5E",x"66",x"5D",x"54",x"0A",x"0A",x"00",x"00",x"00",x"00",x"00", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"13",x"13",x"13",x"13",x"13",x"12",x"12",x"12",x"12",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"13",x"54",x"55",x"5E",x"5E",x"66",x"66",x"5E",x"0B",x"0A",x"00",x"00",x"0A",x"0A",x"0A",x"0A",x"0A",x"0B",x"0B",x"0B",x"0B",x"0C",x"14",x"5D",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"56",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"5E",x"67",x"66",x"66",x"66",x"66",x"66",x"66",x"66",x"66",x"67",x"A7",x"67",x"66",x"66",x"66",x"5E",x"55",x"14",x"14",x"55",x"5D",x"66",x"65",x"5C",x"0A",x"0A",x"0A",x"00",x"00",x"00",x"00", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"12",x"12",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"13",x"14",x"55",x"5E",x"5E",x"66",x"66",x"5E",x"0B",x"0A",x"00",x"00",x"0A",x"0A",x"0A",x"0A",x"0A",x"0B",x"0B",x"0B",x"0B",x"14",x"14",x"55",x"5D",x"5E",x"5E",x"5E",x"5E",x"5F",x"56",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"5E",x"66",x"66",x"66",x"66",x"66",x"66",x"66",x"66",x"66",x"67",x"A7",x"66",x"66",x"66",x"66",x"5E",x"5D",x"0C",x"14",x"15",x"5D",x"66",x"65",x"5D",x"0A",x"0A",x"0A",x"00",x"00",x"00",x"00", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"0C",x"0C",x"0B",x"13",x"0B",x"0B",x"0B",x"13",x"13",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0B",x"14",x"55",x"5E",x"5E",x"5E",x"66",x"66",x"0B",x"0A",x"00",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0B",x"0B",x"0B",x"14",x"14",x"55",x"5D",x"5D",x"5E",x"5E",x"5E",x"5E",x"5F",x"5F",x"56",x"0D",x"0D",x"0D",x"01",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"5E",x"5E",x"67",x"66",x"66",x"66",x"66",x"66",x"66",x"66",x"66",x"66",x"66",x"66",x"66",x"66",x"5E",x"5D",x"55",x"14",x"55",x"5D",x"5D",x"66",x"5D",x"53",x"0A",x"0A",x"00",x"00",x"00",x"00", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"4C",x"0C",x"0C",x"0C",x"0C",x"0B",x"0B",x"0B",x"13",x"0B",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0B",x"54",x"55",x"5E",x"5E",x"5E",x"66",x"66",x"0B",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0B",x"0B",x"0B",x"14",x"14",x"54",x"55",x"5D",x"5E",x"5E",x"5E",x"5E",x"5E",x"5F",x"5E",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"5E",x"5E",x"66",x"5E",x"66",x"66",x"66",x"66",x"66",x"66",x"66",x"66",x"66",x"66",x"66",x"66",x"5E",x"5D",x"5D",x"14",x"15",x"55",x"5D",x"66",x"65",x"54",x"0A",x"0A",x"00",x"00",x"00",x"00", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"55",x"55",x"55",x"15",x"14",x"14",x"0C",x"0B",x"0B",x"0B",x"0B",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"13",x"54",x"55",x"5E",x"5E",x"5E",x"66",x"66",x"0C",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0B",x"0B",x"13",x"14",x"14",x"14",x"55",x"5D",x"5D",x"5E",x"5E",x"5E",x"5E",x"5F",x"5F",x"56",x"0D",x"0C",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"5E",x"5E",x"66",x"5E",x"5E",x"5E",x"66",x"66",x"66",x"66",x"66",x"66",x"A7",x"66",x"66",x"66",x"66",x"5D",x"5D",x"14",x"15",x"14",x"5E",x"66",x"66",x"5D",x"0A",x"0A",x"00",x"00",x"00",x"00", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"4D",x"55",x"55",x"55",x"55",x"55",x"15",x"0C",x"0B",x"0B",x"0B",x"0B",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"13",x"55",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"54",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0B",x"0B",x"14",x"14",x"14",x"14",x"55",x"55",x"5D",x"5E",x"5E",x"5E",x"5E",x"5E",x"5F",x"5E",x"0D",x"0C",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"56",x"5E",x"5E",x"5E",x"5E",x"5E",x"66",x"66",x"66",x"66",x"66",x"66",x"A7",x"66",x"66",x"66",x"66",x"5E",x"5D",x"14",x"5D",x"14",x"66",x"66",x"65",x"65",x"0B",x"0A",x"0A",x"00",x"00",x"00", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"0D",x"0D",x"56",x"55",x"55",x"56",x"55",x"55",x"0C",x"0C",x"0B",x"0B",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"13",x"55",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"54",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0B",x"14",x"54",x"14",x"15",x"55",x"55",x"55",x"5D",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"55",x"0C",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0C",x"55",x"5D",x"5E",x"5E",x"5E",x"5E",x"66",x"66",x"66",x"66",x"66",x"A6",x"AF",x"66",x"66",x"66",x"66",x"66",x"5D",x"14",x"55",x"14",x"66",x"66",x"65",x"65",x"13",x"0A",x"0A",x"00",x"00",x"00", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"0D",x"0D",x"0D",x"0D",x"16",x"56",x"56",x"56",x"56",x"55",x"0C",x"0B",x"0B",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"13",x"55",x"5E",x"5E",x"5E",x"5E",x"5E",x"66",x"5D",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0B",x"0B",x"54",x"54",x"55",x"55",x"55",x"55",x"5D",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"0D",x"0C",x"0C",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0C",x"55",x"55",x"5E",x"5E",x"5E",x"5E",x"5E",x"66",x"66",x"66",x"66",x"A7",x"AF",x"66",x"66",x"66",x"66",x"66",x"5D",x"14",x"14",x"55",x"66",x"66",x"66",x"65",x"53",x"0A",x"0A",x"00",x"00",x"00", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"0D",x"0D",x"0D",x"0D",x"0E",x"0E",x"16",x"56",x"56",x"55",x"55",x"0C",x"0B",x"0B",x"0A",x"0A",x"0A",x"0A",x"0A",x"0B",x"55",x"5E",x"5E",x"5E",x"5E",x"5E",x"67",x"5D",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0B",x"0B",x"54",x"54",x"55",x"55",x"55",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"55",x"0D",x"0C",x"0C",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0C",x"55",x"55",x"5D",x"5D",x"5E",x"5E",x"5E",x"66",x"66",x"66",x"66",x"A7",x"A7",x"66",x"66",x"66",x"66",x"66",x"5D",x"14",x"14",x"5D",x"66",x"66",x"66",x"65",x"53",x"0A",x"0A",x"00",x"00",x"00", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"0D",x"0D",x"0D",x"0D",x"0E",x"0E",x"0E",x"16",x"16",x"56",x"56",x"55",x"0C",x"0B",x"0B",x"0B",x"0A",x"0A",x"0A",x"0B",x"55",x"5E",x"5E",x"5E",x"5E",x"5E",x"67",x"5E",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0B",x"0B",x"54",x"55",x"55",x"5D",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"66",x"5E",x"5E",x"5E",x"5E",x"15",x"0C",x"0C",x"0C",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0C",x"0C",x"0C",x"55",x"15",x"55",x"5D",x"5E",x"5E",x"5E",x"5E",x"66",x"66",x"66",x"A6",x"A7",x"66",x"66",x"66",x"66",x"66",x"5D",x"14",x"55",x"66",x"66",x"66",x"A6",x"5D",x"53",x"0A",x"0A",x"00",x"00",x"00", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0E",x"0E",x"4E",x"4E",x"55",x"55",x"4D",x"0C",x"0B",x"0B",x"0A",x"0B",x"0B",x"54",x"5D",x"5E",x"67",x"5E",x"5E",x"67",x"5E",x"0B",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0B",x"0B",x"14",x"55",x"5D",x"5D",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"55",x"0D",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"15",x"55",x"55",x"5D",x"5E",x"5E",x"5E",x"5E",x"66",x"66",x"66",x"A6",x"A7",x"66",x"66",x"66",x"5E",x"5D",x"5D",x"14",x"5E",x"66",x"66",x"66",x"65",x"5D",x"5C",x"0A",x"0A",x"00",x"00",x"00", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"0D",x"0D",x"0D",x"0D",x"0D",x"0D",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"4D",x"0D",x"0C",x"0C",x"0B",x"0B",x"0B",x"0B",x"54",x"5D",x"5E",x"5E",x"5E",x"5E",x"66",x"5D",x"13",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0B",x"0B",x"14",x"14",x"55",x"5D",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"56",x"15",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"14",x"55",x"55",x"5D",x"5E",x"5E",x"5E",x"5E",x"66",x"66",x"66",x"A6",x"A7",x"66",x"66",x"66",x"5E",x"5D",x"5D",x"14",x"5E",x"66",x"66",x"66",x"65",x"5D",x"5D",x"0A",x"0A",x"00",x"00",x"00", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"0D",x"0D",x"4D",x"4D",x"0D",x"0D",x"0E",x"0E",x"0E",x"0E",x"0D",x"0D",x"0D",x"0D",x"0D",x"0C",x"0B",x"0B",x"0B",x"0B",x"54",x"5E",x"5E",x"5E",x"5E",x"5E",x"66",x"5D",x"13",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0B",x"0B",x"14",x"15",x"55",x"5D",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"56",x"0D",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0B",x"0C",x"0C",x"14",x"55",x"55",x"5D",x"5E",x"5E",x"5E",x"5E",x"66",x"66",x"66",x"66",x"A7",x"66",x"66",x"66",x"5E",x"5D",x"5D",x"14",x"5E",x"66",x"66",x"66",x"66",x"65",x"5D",x"0A",x"0A",x"00",x"00",x"00", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"0D",x"0D",x"4E",x"4E",x"4E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0D",x"0D",x"0D",x"4D",x"55",x"0B",x"0B",x"0B",x"0C",x"55",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5D",x"0B",x"0A",x"0A",x"0A",x"0A",x"0A",x"0B",x"0B",x"13",x"14",x"55",x"5D",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"55",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0B",x"0B",x"0C",x"0C",x"55",x"55",x"5D",x"5E",x"5E",x"5E",x"5E",x"5E",x"66",x"66",x"66",x"66",x"66",x"66",x"66",x"5E",x"5D",x"55",x"14",x"5E",x"66",x"66",x"66",x"66",x"66",x"5D",x"0B",x"0A",x"00",x"00",x"00", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"0E",x"4E",x"4E",x"4E",x"4E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0D",x"4D",x"55",x"55",x"14",x"0B",x"0B",x"55",x"5D",x"5E",x"5E",x"5E",x"5E",x"5E",x"66",x"5D",x"0B",x"0A",x"0A",x"0A",x"0A",x"0A",x"0B",x"0B",x"14",x"54",x"55",x"5D",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5D",x"15",x"0C",x"0B",x"0B",x"0B",x"0B",x"0C",x"0B",x"0B",x"0B",x"0C",x"14",x"55",x"55",x"5D",x"5D",x"5E",x"5E",x"5E",x"5E",x"5E",x"66",x"66",x"66",x"66",x"66",x"5E",x"5E",x"5D",x"14",x"14",x"5E",x"66",x"66",x"66",x"66",x"66",x"5D",x"13",x"0A",x"00",x"00",x"00", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"0E",x"0E",x"4E",x"4E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0D",x"0D",x"4D",x"55",x"54",x"14",x"54",x"5D",x"5E",x"5E",x"5E",x"5E",x"5F",x"67",x"66",x"5D",x"14",x"0A",x"0A",x"0A",x"0A",x"0A",x"0B",x"0B",x"14",x"54",x"55",x"5D",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"55",x"0C",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0B",x"0C",x"14",x"54",x"55",x"5D",x"5D",x"5D",x"5E",x"5E",x"5E",x"5E",x"5E",x"66",x"66",x"5E",x"66",x"5E",x"5E",x"5E",x"14",x"55",x"5E",x"66",x"5D",x"5D",x"66",x"A6",x"65",x"54",x"0A",x"0A",x"00",x"00", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"0E",x"0E",x"0E",x"0E",x"0E",x"16",x"16",x"16",x"0E",x"0E",x"0E",x"0E",x"0D",x"0D",x"0D",x"4D",x"0C",x"55",x"5D",x"5E",x"5E",x"5E",x"5E",x"5E",x"5F",x"67",x"66",x"5E",x"54",x"0A",x"0A",x"0A",x"0A",x"0A",x"0B",x"0B",x"14",x"55",x"55",x"5D",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5D",x"14",x"0B",x"0A",x"0B",x"0B",x"0A",x"0A",x"0B",x"0B",x"0B",x"14",x"54",x"55",x"5D",x"5D",x"5D",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"66",x"5E",x"66",x"5E",x"5E",x"5E",x"14",x"55",x"5E",x"5E",x"5D",x"5D",x"65",x"A6",x"66",x"5C",x"0A",x"0A",x"00",x"00", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"0E",x"0E",x"0E",x"0E",x"0E",x"16",x"16",x"16",x"16",x"56",x"56",x"0E",x"0D",x"0D",x"0C",x"0C",x"0C",x"55",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"67",x"67",x"5E",x"5E",x"5D",x"0B",x"0A",x"0A",x"0A",x"0A",x"0B",x"0B",x"14",x"55",x"55",x"5D",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5D",x"54",x"0B",x"0A",x"0A",x"0A",x"0A",x"0B",x"0B",x"0B",x"0B",x"54",x"14",x"14",x"55",x"55",x"5D",x"5D",x"5E",x"5E",x"5E",x"5E",x"5E",x"66",x"5E",x"66",x"5E",x"5E",x"5E",x"14",x"5D",x"5D",x"5D",x"54",x"54",x"5D",x"66",x"66",x"5D",x"0A",x"0A",x"0A",x"00", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"0D",x"0E",x"0E",x"16",x"16",x"16",x"16",x"56",x"56",x"57",x"5F",x"56",x"0D",x"0C",x"01",x"0C",x"0C",x"5D",x"5E",x"5E",x"5D",x"5E",x"5E",x"5E",x"67",x"67",x"67",x"5E",x"5D",x"54",x"0A",x"0A",x"0A",x"0A",x"0B",x"0B",x"14",x"55",x"55",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5D",x"5D",x"54",x"0B",x"0A",x"0A",x"0A",x"0A",x"0A",x"0B",x"0B",x"0B",x"14",x"54",x"54",x"55",x"55",x"55",x"5D",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5D",x"55",x"5D",x"66",x"54",x"13",x"13",x"5D",x"A6",x"A6",x"65",x"5B",x"0A",x"0A",x"00", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"0D",x"0D",x"0E",x"0E",x"16",x"16",x"16",x"16",x"56",x"57",x"57",x"56",x"0D",x"0C",x"01",x"0C",x"0C",x"5E",x"5E",x"5E",x"5D",x"5D",x"5E",x"5E",x"67",x"67",x"67",x"5E",x"5E",x"5D",x"0B",x"0A",x"0A",x"0A",x"0B",x"0B",x"14",x"55",x"55",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5D",x"5D",x"13",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0B",x"0B",x"13",x"54",x"54",x"55",x"55",x"55",x"5D",x"5D",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5D",x"55",x"5D",x"66",x"54",x"0B",x"0B",x"5C",x"A6",x"66",x"5D",x"53",x"0A",x"0A",x"00", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"0D",x"0D",x"0D",x"0E",x"16",x"16",x"16",x"16",x"56",x"56",x"56",x"55",x"0C",x"01",x"01",x"0B",x"0C",x"5E",x"5E",x"5E",x"5D",x"55",x"5E",x"67",x"67",x"67",x"67",x"5E",x"5E",x"5D",x"54",x"0A",x"0A",x"0A",x"0B",x"0B",x"14",x"54",x"55",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5D",x"5D",x"0B",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0B",x"0B",x"0B",x"14",x"54",x"54",x"55",x"55",x"55",x"5D",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"55",x"55",x"5D",x"5D",x"0B",x"0A",x"0A",x"5C",x"65",x"5E",x"5C",x"52",x"4A",x"0A",x"0A", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--        x"0D",x"0D",x"0D",x"0D",x"0D",x"16",x"16",x"16",x"56",x"56",x"56",x"0D",x"0C",x"0C",x"01",x"0B",x"0C",x"55",x"5D",x"5E",x"5E",x"55",x"5E",x"67",x"67",x"5E",x"67",x"5E",x"5E",x"66",x"5D",x"0A",x"0A",x"0A",x"0B",x"0B",x"14",x"54",x"55",x"5D",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5D",x"5D",x"0B",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0B",x"0B",x"0B",x"14",x"54",x"54",x"55",x"55",x"55",x"5D",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"5E",x"15",x"5D",x"5E",x"5D",x"0B",x"0A",x"0A",x"5C",x"65",x"5D",x"54",x"53",x"52",x"52",x"0A", x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
--    others=>x"00");
    
            
    begin
    -- Process to control the memory access
    process(clk)
    begin
        if rising_edge(clk) then    -- Memory writing        
            if we = '1' then
                RAM(TO_INTEGER(UNSIGNED(address))) <= data_in; 
            end if;
            -- Synchronous memory read (Block RAM)
            data_out <= RAM(TO_INTEGER(UNSIGNED(address)));
        end if;   
    end process;
    
end BLOCK_RAM;