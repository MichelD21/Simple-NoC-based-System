-- ######################################################
-- #          < STORM SoC by Stephan Nolting >          #
-- # ************************************************** #
-- #             Internal Memory Component              #
-- # ************************************************** #
-- # Last modified: 04.03.2012                          #
-- ######################################################

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;


entity MEMORY is
	generic	(
				MEM_SIZE      : natural := 256;  -- memory cells
				LOG2_MEM_SIZE : natural := 8;    -- log2(memory cells)
				OUTPUT_GATE   : boolean := FALSE -- output and-gate, might be necessary for some bus systems
			);
	port	(
				-- Wishbone Bus --
				WB_CLK_I      : in  STD_LOGIC; -- memory master clock
				WB_RST_I      : in  STD_LOGIC; -- high active sync reset
				WB_CTI_I      : in  STD_LOGIC_VECTOR(02 downto 0); -- cycle indentifier
				WB_TGC_I      : in  STD_LOGIC_VECTOR(06 downto 0); -- cycle tag
				WB_ADR_I      : in  STD_LOGIC_VECTOR(LOG2_MEM_SIZE-1 downto 0); -- adr in
				WB_DATA_I     : in  STD_LOGIC_VECTOR(31 downto 0); -- write data
				WB_DATA_O     : out STD_LOGIC_VECTOR(31 downto 0); -- read data
				WB_SEL_I      : in  STD_LOGIC_VECTOR(03 downto 0); -- data quantity
				WB_WE_I       : in  STD_LOGIC; -- write enable
				WB_STB_I      : in  STD_LOGIC; -- valid cycle
				WB_ACK_O      : out STD_LOGIC; -- acknowledge
				WB_HALT_O     : out STD_LOGIC; -- throttle master
				WB_ERR_O      : out STD_LOGIC  -- abnormal cycle termination
			);
end MEMORY;

architecture Behavioral of MEMORY is

	--- Buffer ---
	signal WB_ACK_O_INT : STD_LOGIC;
	signal WB_DATA_INT  : STD_LOGIC_VECTOR(31 downto 0);

	--- Memory Type ---
	type MEM_FILE_TYPE is array (0 to MEM_SIZE - 1) of STD_LOGIC_VECTOR(31 downto 0);

	--- INIT MEMORY IMAGE ---
	------------------------------------------------------
	signal MEM_FILE : MEM_FILE_TYPE :=
	(
		000000 => x"E10F1000",
000001 => x"E3C11080",
000002 => x"E121F001",
000003 => x"EB000000",
000004 => x"EAFFFFFE",
000005 => x"E3E03A01",
000006 => x"E5132FDB",
000007 => x"E3A02B01",
000008 => x"E92D41F0",
000009 => x"E5032FDF",
000010 => x"E3A06000",
000011 => x"E59F8228",
000012 => x"E1A07006",
000013 => x"E087E008",
000014 => x"E3A0C000",
000015 => x"E3865C06",
000016 => x"E3864B01",
000017 => x"E3E02A01",
000018 => x"E5123FDB",
000019 => x"E3130B01",
000020 => x"0AFFFFFC",
000021 => x"E3A03C06",
000022 => x"E3A02B01",
000023 => x"E3E01A01",
000024 => x"E2833003",
000025 => x"E2822003",
000026 => x"E5013FDF",
000027 => x"E5012FDF",
000028 => x"E5113FDB",
000029 => x"E3130B01",
000030 => x"1A000003",
000031 => x"E1A02001",
000032 => x"E5123FDB",
000033 => x"E3130B01",
000034 => x"0AFFFFFC",
000035 => x"E1A03A85",
000036 => x"E1A02A84",
000037 => x"E3E01A01",
000038 => x"E1A03AA3",
000039 => x"E1A02AA2",
000040 => x"E5013FDF",
000041 => x"E5012FDF",
000042 => x"E5113FDB",
000043 => x"E3130B01",
000044 => x"1A000003",
000045 => x"E1A02001",
000046 => x"E5123FDB",
000047 => x"E3130B01",
000048 => x"0AFFFFFC",
000049 => x"E38C3C06",
000050 => x"E38C2B01",
000051 => x"E1A03A83",
000052 => x"E1A02A82",
000053 => x"E3E01A01",
000054 => x"E1A03AA3",
000055 => x"E1A02AA2",
000056 => x"E5013FDF",
000057 => x"E5012FDF",
000058 => x"E5113FDB",
000059 => x"E3130B01",
000060 => x"E5DE0000",
000061 => x"1A000003",
000062 => x"E1A02001",
000063 => x"E5123FDB",
000064 => x"E3130B01",
000065 => x"0AFFFFFC",
000066 => x"E28CC001",
000067 => x"E3E02A01",
000068 => x"E3801B01",
000069 => x"E3803C07",
000070 => x"E35C0032",
000071 => x"E5023FDF",
000072 => x"E28EE001",
000073 => x"E5021FDF",
000074 => x"1AFFFFC5",
000075 => x"E2866001",
000076 => x"E3560032",
000077 => x"E2877032",
000078 => x"1AFFFFBD",
000079 => x"E3A07000",
000080 => x"E3A06064",
000081 => x"E087E008",
000082 => x"E3A0C000",
000083 => x"E3865C06",
000084 => x"E3864B01",
000085 => x"E3E02A01",
000086 => x"E5123FDB",
000087 => x"E3130B01",
000088 => x"0AFFFFFC",
000089 => x"E3A03C06",
000090 => x"E3A02B01",
000091 => x"E3E01A01",
000092 => x"E2833003",
000093 => x"E2822003",
000094 => x"E5013FDF",
000095 => x"E5012FDF",
000096 => x"E5113FDB",
000097 => x"E3130B01",
000098 => x"1A000003",
000099 => x"E1A02001",
000100 => x"E5123FDB",
000101 => x"E3130B01",
000102 => x"0AFFFFFC",
000103 => x"E1A03A85",
000104 => x"E1A02A84",
000105 => x"E3E01A01",
000106 => x"E1A03AA3",
000107 => x"E1A02AA2",
000108 => x"E5013FDF",
000109 => x"E5012FDF",
000110 => x"E5113FDB",
000111 => x"E3130B01",
000112 => x"1A000003",
000113 => x"E1A02001",
000114 => x"E5123FDB",
000115 => x"E3130B01",
000116 => x"0AFFFFFC",
000117 => x"E38C3C06",
000118 => x"E38C2B01",
000119 => x"E1A03A83",
000120 => x"E1A02A82",
000121 => x"E3E01A01",
000122 => x"E1A03AA3",
000123 => x"E1A02AA2",
000124 => x"E5013FDF",
000125 => x"E5012FDF",
000126 => x"E5113FDB",
000127 => x"E3130B01",
000128 => x"E5DE0000",
000129 => x"1A000003",
000130 => x"E1A02001",
000131 => x"E5123FDB",
000132 => x"E3130B01",
000133 => x"0AFFFFFC",
000134 => x"E28CC001",
000135 => x"E3E02A01",
000136 => x"E3801B01",
000137 => x"E3803C07",
000138 => x"E35C0032",
000139 => x"E5023FDF",
000140 => x"E28EE001",
000141 => x"E5021FDF",
000142 => x"1AFFFFC5",
000143 => x"E3A03D27",
000144 => x"E2877032",
000145 => x"E2833004",
000146 => x"E1570003",
000147 => x"E2866001",
000148 => x"1AFFFFBB",
000149 => x"E3A00000",
000150 => x"E8BD81F0",
000151 => x"00000360",
000152 => x"00000000",
000153 => x"00000000",
000154 => x"00000000",
000155 => x"00000000",
000156 => x"00000000",
000157 => x"00000000",
000158 => x"00000000",
000159 => x"00000000",
000160 => x"00000000",
000161 => x"00000000",
000162 => x"00000000",
000163 => x"00000000",
000164 => x"00000000",
000165 => x"00000000",
000166 => x"00000000",
000167 => x"00000000",
000168 => x"00000000",
000169 => x"00000000",
000170 => x"00000000",
000171 => x"00000000",
000172 => x"00000000",
000173 => x"00000000",
000174 => x"00000000",
000175 => x"00000000",
000176 => x"00000000",
000177 => x"00000000",
000178 => x"00000000",
000179 => x"00000000",
000180 => x"00000000",
000181 => x"00000000",
000182 => x"00000000",
000183 => x"00000000",
000184 => x"00000000",
000185 => x"00000000",
000186 => x"00000000",
000187 => x"00000000",
000188 => x"00000000",
000189 => x"00000000",
000190 => x"00000000",
000191 => x"00000000",
000192 => x"00000000",
000193 => x"00000000",
000194 => x"00000000",
000195 => x"00000000",
000196 => x"00000000",
000197 => x"00000000",
000198 => x"00000000",
000199 => x"00000000",
000200 => x"00000000",
000201 => x"00000000",
000202 => x"00000000",
000203 => x"00000000",
000204 => x"00000000",
000205 => x"00000000",
000206 => x"00000000",
000207 => x"00000000",
000208 => x"00000000",
000209 => x"00000000",
000210 => x"00000000",
000211 => x"00000000",
000212 => x"00000000",
000213 => x"00000000",
000214 => x"00000000",
000215 => x"00000000",
000216 => x"54540A00",
000217 => x"00000000",
000218 => x"00000A0A",
000219 => x"0A0A0000",
000220 => x"0A0A0A0B",
000221 => x"0B0B0B0B",
000222 => x"0B0A0A00",
000223 => x"0A0A0A0A",
000224 => x"0A0A0B4B",
000225 => x"0A000000",
000226 => x"00000000",
000227 => x"0000000A",
000228 => x"0A0B540C",
000229 => x"0A000000",
000230 => x"0A4C554D",
000231 => x"0A555554",
000232 => x"0A0A545C",
000233 => x"4C0B4C55",
000234 => x"55550C0B",
000235 => x"0A54540B",
000236 => x"0A0A0B0B",
000237 => x"5D540A00",
000238 => x"545C540A",
000239 => x"5C540000",
000240 => x"000A0A0C",
000241 => x"4B0B0A00",
000242 => x"00000B4D",
000243 => x"0B010B0B",
000244 => x"0B4C0A54",
000245 => x"4A0A4C0C",
000246 => x"0B0B4B0B",
000247 => x"55010B0B",
000248 => x"4B540A0A",
000249 => x"544C0B0A",
000250 => x"0B004C0A",
000251 => x"0A4D4A0B",
000252 => x"0000000A",
000253 => x"0A0C0A0A",
000254 => x"0A0A0000",
000255 => x"0A54F69D",
000256 => x"55FFF755",
000257 => x"004BF6F6",
000258 => x"0B559DF6",
000259 => x"F6F6074B",
000260 => x"0A07F654",
000261 => x"0A0B1455",
000262 => x"F607550A",
000263 => x"4CF6A54E",
000264 => x"F6070000",
000265 => x"00000A0B",
000266 => x"000A0A0A",
000267 => x"0A000A55",
000268 => x"F6AF4CFF",
000269 => x"A45E004B",
000270 => x"F6F60B55",
000271 => x"9DFFF6F6",
000272 => x"F60A0B07",
000273 => x"F6540A0B",
000274 => x"0C55F607",
000275 => x"9E0A4CFF",
000276 => x"A54EF6EE",
000277 => x"00000000",
000278 => x"0A0B000A",
000279 => x"4A0A0A00",
000280 => x"000AF6F6",
000281 => x"0AF60B01",
000282 => x"0A43F6F6",
000283 => x"4C559DF6",
000284 => x"A5F6FF9C",
000285 => x"0C07F654",
000286 => x"0A0B0D4D",
000287 => x"F6074C00",
000288 => x"4BFF9D56",
000289 => x"F6AE0000",
000290 => x"0000000A",
000291 => x"000A0A0A",
000292 => x"0A000A0A",
000293 => x"07FFFFF7",
000294 => x"0C0B0CAE",
000295 => x"F6F60754",
000296 => x"A5FFAE54",
000297 => x"F6AD4D08",
000298 => x"F6550A0C",
000299 => x"0D4BF6F6",
000300 => x"4B0C4BFF",
000301 => x"5C56FF08",
000302 => x"00000000",
000303 => x"0000000A",
000304 => x"0B0B0A00",
000305 => x"9D0AAEF6",
000306 => x"FF9C0B14",
000307 => x"0D07A4FF",
000308 => x"0755A5F6",
000309 => x"5C07F654",
000310 => x"0E08F655",
000311 => x"0A15565C",
000312 => x"F7F6544D",
000313 => x"4BFF5C56",
000314 => x"F6F70A00",
000315 => x"00000000",
000316 => x"000A0B4C",
000317 => x"0B0A5D53",
000318 => x"5DF6FF53",
000319 => x"0B150DF6",
000320 => x"5BFF0854",
000321 => x"9DF6EFF6",
000322 => x"F64B0E08",
000323 => x"F6550A55",
000324 => x"569DA5F6",
000325 => x"5C554CFF",
000326 => x"5C4EF6F7",
000327 => x"00000000",
000328 => x"00000A0B",
000329 => x"0C540C54",
000330 => x"00000BF6",
000331 => x"F64C0C15",
000332 => x"57084AF6",
000333 => x"085E9CFF",
000334 => x"08FF084C",
000335 => x"0EF6F655",
000336 => x"0A5D56F6",
000337 => x"9BF6AE56",
000338 => x"4CFF9D4D",
000339 => x"F6F70A0A",
000340 => x"0A0A0A00",
000341 => x"0A0B0C55",
000342 => x"0C0B0A00",
000343 => x"5DFFF60A",
000344 => x"0C5E1508",
000345 => x"0A08F654",
000346 => x"5CFF0808",
000347 => x"08530EF6",
000348 => x"F6550A56",
000349 => x"4CF653F6",
000350 => x"F7544CF6",
000351 => x"AE4EF6F7",
000352 => x"0A0A0A0A",
000353 => x"0A0A0C0C",
000354 => x"0C550C0B",
000355 => x"0A0AF6F6",
000356 => x"F69D0D15",
000357 => x"15F607F6",
000358 => x"F6AF5CF6",
000359 => x"9D0AF6F6",
000360 => x"5607FF56",
000361 => x"0B0C0BF6",
000362 => x"07F6080B",
000363 => x"01F65C57",
000364 => x"F6F70A0A",
000365 => x"0A0A0A0A",
000366 => x"0C0C0C55",
000367 => x"0C0B0A0A",
000368 => x"08F6F6A6",
000369 => x"0D1E15F6",
000370 => x"08FFF65E",
000371 => x"9DF69D0B",
000372 => x"F6F65608",
000373 => x"F6560B0C",
000374 => x"0AF608F6",
000375 => x"080B0CF6",
000376 => x"9D57F6F7",
000377 => x"0A0A0A0A",
000378 => x"0A0A155E",
000379 => x"5E0C0C0B",
000380 => x"0B55F6F6",
000381 => x"53F60C16",
000382 => x"55FF54F7",
000383 => x"FF5E5CFF",
000384 => x"F653F607",
000385 => x"5F07F64C",
000386 => x"54015DF6",
000387 => x"53F6F65C",
000388 => x"4CF6A456",
000389 => x"F6F70A0A",
000390 => x"0A0A0A0A",
000391 => x"151E550C",
000392 => x"0C0B0B15",
000393 => x"F6F654F6",
000394 => x"A7160DF6",
000395 => x"545CF656",
000396 => x"9DF6A507",
000397 => x"F6070D07",
000398 => x"F60A0A55",
000399 => x"A6F654F6",
000400 => x"F6A54DF6",
000401 => x"074CF6AD",
000402 => x"0A0A0A0A",
000403 => x"0A0A1455",
000404 => x"0D0C0C0B",
000405 => x"0C55F6A5",
000406 => x"5E08AE56",
000407 => x"EFF64D0B",
000408 => x"F65F5DF6",
000409 => x"F6F6F6B7",
000410 => x"AF07F6F6",
000411 => x"F656F6F6",
000412 => x"5607F6EE",
000413 => x"5508F6F6",
000414 => x"07530A0A",
000415 => x"0A0C0A0A",
000416 => x"0C675655",
000417 => x"5514554C",
000418 => x"074B5607",
000419 => x"EE015C08",
000420 => x"550B075E",
000421 => x"5DF608F6",
000422 => x"EF1CF608",
000423 => x"08080855",
000424 => x"9B0855A5",
000425 => x"08074D4B",
000426 => x"08084B54",
000427 => x"0B0B0B0B",
000428 => x"0A0A145E",
000429 => x"5E561515",
000430 => x"67550A0C",
000431 => x"160B0B0C",
000432 => x"0C0BA715",
000433 => x"0A56010B",
000434 => x"0A0A4C1E",
000435 => x"B70B0A5C",
000436 => x"0A560B0A",
000437 => x"4D0B0A0A",
000438 => x"0C540B0B",
000439 => x"540B0B0B",
000440 => x"0B0B0A0A",
000441 => x"0C155E5E",
000442 => x"1E676F6F",
000443 => x"67B71615",
000444 => x"15151516",
000445 => x"1515162F",
000446 => x"2F272727",
000447 => x"27272F1E",
000448 => x"1E1E1E15",
000449 => x"14151515",
000450 => x"15151515",
000451 => x"1455151E",
000452 => x"1514140C",
000453 => x"0B0A0C15",
000454 => x"5E5E1E67",
000455 => x"6F6F676F",
000456 => x"16151515",
000457 => x"15151515",
000458 => x"1E2F2F27",
000459 => x"6767272F",
000460 => x"2F1F1E1E",
000461 => x"1F151E15",
000462 => x"15151515",
000463 => x"16150C14",
000464 => x"151E1615",
000465 => x"150C0B0A",
000466 => x"1515151E",
000467 => x"1E676F6F",
000468 => x"271E1615",
000469 => x"15151515",
000470 => x"16161E6F",
000471 => x"2F2F6F6F",
000472 => x"6F6F6F6F",
000473 => x"B766671E",
000474 => x"6F6F1E15",
000475 => x"151E5F16",
000476 => x"15151515",
000477 => x"150C140C",
000478 => x"0B0A1515",
000479 => x"151E1E27",
000480 => x"6F6F1E1E",
000481 => x"16151515",
000482 => x"15161E1E",
000483 => x"1F6F2F6F",
000484 => x"6FB7B76F",
000485 => x"6FAFB7B7",
000486 => x"B71E2727",
000487 => x"6715151E",
000488 => x"1F161515",
000489 => x"15151555",
000490 => x"14140B0A",
000491 => x"1515551E",
000492 => x"1F1F6F6F",
000493 => x"1F1F1E15",
000494 => x"1515151E",
000495 => x"1E1E272F",
000496 => x"77BFEF5D",
000497 => x"EEF6F6B6",
000498 => x"AFAEF66F",
000499 => x"272F6F1E",
000500 => x"1E1E6F27",
000501 => x"1E165656",
000502 => x"0E564D15",
000503 => x"0C0A1515",
000504 => x"551E1F1F",
000505 => x"6F6F1F1F",
000506 => x"1E151515",
000507 => x"151E1E1E",
000508 => x"272F77BF",
000509 => x"EF5DEEF6",
000510 => x"F6B6AFAE",
000511 => x"F66F272F",
000512 => x"6F1E1E1E",
000513 => x"6F271E16",
000514 => x"56560E56",
000515 => x"4D150C0A",
000516 => x"150C0D16",
000517 => x"161F2F6F",
000518 => x"1F1F1E16",
000519 => x"161E1F1F",
000520 => x"2727276F",
000521 => x"6FF6F65C",
000522 => x"07EFB7B7",
000523 => x"A5F6F6B7",
000524 => x"6F6F6F27",
000525 => x"272F7727",
000526 => x"1F1E0E4E",
000527 => x"4E4D4E15",
000528 => x"0C0B1555",
000529 => x"4D56561E",
000530 => x"2F2F2727",
000531 => x"271E1E1F",
000532 => x"1F272727",
000533 => x"2F776FF6",
000534 => x"F608F6AF",
000535 => x"67AFF6F6",
000536 => x"F6AF6F6F",
000537 => x"6F6F2F6F",
000538 => x"77271E1F",
000539 => x"0E0E0E4E",
000540 => x"5515140C",
000541 => x"154D4E4E",
000542 => x"4E5E2F2F",
000543 => x"271F2727",
000544 => x"271E2727",
000545 => x"27272F6F",
000546 => x"66F6F6F6",
000547 => x"B7675F67",
000548 => x"EFF6F6AF",
000549 => x"67672F77",
000550 => x"6F777727",
000551 => x"1E1F0E4E",
000552 => x"0E0D1515",
000553 => x"140C1E0D",
000554 => x"4D4D4D56",
000555 => x"2F272727",
000556 => x"27272727",
000557 => x"27272727",
000558 => x"2767555D",
000559 => x"A55D551F",
000560 => x"1F5F56AF",
000561 => x"EF55561E",
000562 => x"77777777",
000563 => x"7727275F",
000564 => x"0D0D0D15",
000565 => x"67151415",
000566 => x"1E0D4D4D",
000567 => x"4D152727",
000568 => x"27272727",
000569 => x"27672727",
000570 => x"2727275E",
000571 => x"1554544C",
000572 => x"0D1F1F5F",
000573 => x"55A6AF55",
000574 => x"56167777",
000575 => x"77777727",
000576 => x"675F0D0D",
000577 => x"0D155E15",
000578 => x"141D1E56",
000579 => x"550D0D56",
000580 => x"671F2727",
000581 => x"6F6F2767",
000582 => x"27272727",
000583 => x"670D0D01",
000584 => x"0C010117",
000585 => x"17570E0C",
000586 => x"4D0D0D56",
000587 => x"6F777777",
000588 => x"772F671E",
000589 => x"014D151E",
000590 => x"5E14141E",
000591 => x"275E560D",
000592 => x"4D0D155F",
000593 => x"2727776F",
000594 => x"2F2F272F",
000595 => x"27675F4D",
000596 => x"0C010C0C",
000597 => x"010D570E",
000598 => x"0C0B0C0C",
000599 => x"0C4D1F77",
000600 => x"2F2F2F67",
000601 => x"1E0D0D0D",
000602 => x"5E1E1515",
000603 => x"141E275E",
000604 => x"560D4D0D",
000605 => x"155F2727",
000606 => x"776F2F2F",
000607 => x"272F2767",
000608 => x"5F4D0C01",
000609 => x"0C0C010D",
000610 => x"570E0C0B",
000611 => x"0C0C0C4D",
000612 => x"1F772F2F",
000613 => x"2F671E0D",
000614 => x"0D0D5E1E",
000615 => x"1515141E",
000616 => x"27272F6F",
000617 => x"67550D0D",
000618 => x"67672F2F",
000619 => x"2F2F6F1E",
000620 => x"56564E0C",
000621 => x"0B0B0B0B",
000622 => x"0B0B0B0A",
000623 => x"0A0A0A0A",
000624 => x"0B0C4E56",
000625 => x"1F6F6715",
000626 => x"0D0D155E",
000627 => x"1E676715",
000628 => x"1E67272F",
000629 => x"2F6F6F15",
000630 => x"4E0D5E77",
000631 => x"2F2F2F2F",
000632 => x"6F56564E",
000633 => x"4E0C0B0C",
000634 => x"0C0C4C4C",
000635 => x"4C0B0B0B",
000636 => x"0B0A0B0C",
000637 => x"4E571F6F",
000638 => x"270D4D0D",
000639 => x"165E1E27",
000640 => x"1655151E",
000641 => x"2F2F2F77",
000642 => x"77670D4D",
000643 => x"0D1E676F",
000644 => x"2F376F16",
000645 => x"0E0E4E0C",
000646 => x"0D0C0D0D",
000647 => x"0C0D0D0D",
000648 => x"0D0D0C0C",
000649 => x"0C0D4E56",
000650 => x"5F6F164D",
000651 => x"4D0D5E1E",
000652 => x"1E151515",
000653 => x"15152F2F",
000654 => x"3777776F",
000655 => x"0D4D0D15",
000656 => x"672F2F37",
000657 => x"6F5F0E0E",
000658 => x"4E0C0D0C",
000659 => x"0D0D0D0D",
000660 => x"0D0D0D0D",
000661 => x"0D0C0C0D",
000662 => x"4E565E67",
000663 => x"164D4D0D",
000664 => x"671E1515",
000665 => x"0D151515",
000666 => x"37373737",
000667 => x"37775F16",
000668 => x"4D0D1577",
000669 => x"77777767",
000670 => x"0D0D0D01",
000671 => x"0101010C",
000672 => x"0C0C0C01",
000673 => x"0D0D0D0D",
000674 => x"0D4D4D0D",
000675 => x"4E564E0D",
000676 => x"0D5E1E1E",
000677 => x"160C0C15",
000678 => x"15153737",
000679 => x"37373737",
000680 => x"671E560D",
000681 => x"0D6F7777",
000682 => x"77670D0D",
000683 => x"0D010101",
000684 => x"010C0101",
000685 => x"0C010D01",
000686 => x"0D0D0D0D",
000687 => x"4D4D0D4E",
000688 => x"4E0D565F",
000689 => x"1E15150C",
000690 => x"0C0C1515",
000691 => x"3777372F",
000692 => x"2F2F776F",
000693 => x"160E4D0D",
000694 => x"6F6F2F6F",
000695 => x"5E4C0C0D",
000696 => x"010C0C01",
000697 => x"01010C0D",
000698 => x"0D0D4D0D",
000699 => x"0C01014D",
000700 => x"4D4E0D16",
000701 => x"67271516",
000702 => x"150C0B0C",
000703 => x"67273737",
000704 => x"7737372F",
000705 => x"3777160E",
000706 => x"0D0D1527",
000707 => x"2F6F670C",
000708 => x"0C4D010C",
000709 => x"0C01010C",
000710 => x"0C0D0D0D",
000711 => x"0D0C0101",
000712 => x"0C0D0D4E",
000713 => x"0D676727",
000714 => x"151E150C",
000715 => x"0C0C6767",
000716 => x"3F7F7737",
000717 => x"372F3777",
000718 => x"5F560D4D",
000719 => x"0D15272F",
000720 => x"670C0101",
000721 => x"010C0C01",
000722 => x"010C0C0D",
000723 => x"0D0D0D01",
000724 => x"010C4C0D",
000725 => x"0D0D566F",
000726 => x"2F271E15",
000727 => x"1E150C55",
000728 => x"6727FB7F",
000729 => x"772F2F27",
000730 => x"2F376F5E",
000731 => x"164D0D0E",
000732 => x"1F6F670C",
000733 => x"0D4D0C0C",
000734 => x"0C010C01",
000735 => x"010D4D0D",
000736 => x"0D010C0C",
000737 => x"0C0D0D0D",
000738 => x"1E6F2F6F",
000739 => x"1F1E165E",
000740 => x"155E6F6F",
000741 => x"3F7F7737",
000742 => x"2F2F2F2F",
000743 => x"6F67164D",
000744 => x"4D0D166F",
000745 => x"670C0D4D",
000746 => x"0C0C0C0C",
000747 => x"0C0C010D",
000748 => x"4D0D0D01",
000749 => x"0C010C0D",
000750 => x"4D0D1E2F",
000751 => x"2F6F1E1F",
000752 => x"155E1567",
000753 => x"6F6FFBFB",
000754 => x"7F777F2F",
000755 => x"372F7F7F",
000756 => x"77564E4E",
000757 => x"0D0C0D4D",
000758 => x"0C4D0D0C",
000759 => x"0D4D0C01",
000760 => x"0C0D0C01",
000761 => x"0C0C0C01",
000762 => x"4C4D0D15",
000763 => x"7737772F",
000764 => x"271E2716",
000765 => x"16672777",
000766 => x"FBFB7F77",
000767 => x"7F2F372F",
000768 => x"7F7F7756",
000769 => x"4E4E0D0C",
000770 => x"0D4D0C4D",
000771 => x"0D0C0D4D",
000772 => x"0C010C0D",
000773 => x"0C010C0C",
000774 => x"0C014C4D",
000775 => x"0D157737",
000776 => x"772F271E",
000777 => x"27161667",
000778 => x"27773F37",
000779 => x"2F27275F",
000780 => x"27277F7F",
000781 => x"7F771E56",
000782 => x"150D0C01",
000783 => x"0C0C0C01",
000784 => x"0101010C",
000785 => x"010C0101",
000786 => x"010C0C01",
000787 => x"0C561E77",
000788 => x"77772F2F",
000789 => x"27675E15",
000790 => x"15151F67",
000791 => x"37372F27",
000792 => x"271E2727",
000793 => x"7F7F7F77",
000794 => x"2656160D",
000795 => x"0C010C01",
000796 => x"0C010C01",
000797 => x"010C0101",
000798 => x"010C0C0D",
000799 => x"0D0C0D56",
000800 => x"1E777777",
000801 => x"2F2F2727",
000802 => x"6715150D",
000803 => x"1E67372F",
000804 => x"2F2F2716",
000805 => x"1E277F7F",
000806 => x"3F777767",
000807 => x"160D0C01",
000808 => x"010C4C0C",
000809 => x"0C0C010C",
000810 => x"0101010C",
000811 => x"010D0D0D",
000812 => x"0D556777",
000813 => x"772F6F6F",
000814 => x"671E675E",
000815 => x"AF0C1567",
000816 => x"372F2727",
000817 => x"271E1F27",
000818 => x"77373777",
000819 => x"7F771E0D",
000820 => x"0C0C0C0C",
000821 => x"0C0C4D0C",
000822 => x"010C0101",
000823 => x"0C0D0D4E",
000824 => x"4D014D0D",
000825 => x"77772F27",
000826 => x"2727671F",
000827 => x"6F5F550C",
000828 => x"0C15376F",
000829 => x"2727271E",
000830 => x"1F677777",
000831 => x"777F7F77",
000832 => x"665F4D4C",
000833 => x"4C0D0C4D",
000834 => x"4D0D0D0D",
000835 => x"0C0C0C0C",
000836 => x"0D0D550D",
000837 => x"555E6F77",
000838 => x"6F27676F",
000839 => x"67676767",
000840 => x"150B0C14",
others => x"F0013007"





);
	------------------------------------------------------

begin

	-- STORM data/instruction memory -----------------------------------------------------------------------
	-- --------------------------------------------------------------------------------------------------------
		MEM_FILE_ACCESS: process(WB_CLK_I)
		begin
			--- Sync Write ---
			if rising_edge(WB_CLK_I) then

				--- Data Read/Write ---
				if (WB_STB_I = '1') then
					if (WB_WE_I = '1') then
						MEM_FILE(to_integer(unsigned(WB_ADR_I))) <= WB_DATA_I;
					end if;
					WB_DATA_INT <= MEM_FILE(to_integer(unsigned(WB_ADR_I)));
				end if;

				--- ACK Control ---
				if (WB_RST_I = '1') then
					WB_ACK_O_INT <= '0';
				elsif (WB_CTI_I = "000") or (WB_CTI_I = "111") then
					WB_ACK_O_INT <= WB_STB_I and (not WB_ACK_O_INT);
				else
					WB_ACK_O_INT <= WB_STB_I;
				end if;

			end if;
		end process MEM_FILE_ACCESS;

		--- Output Gate ---
		WB_DATA_O <= WB_DATA_INT when (OUTPUT_GATE = FALSE) or ((OUTPUT_GATE = TRUE) and (WB_STB_I = '1')) else (others => '0');

		--- ACK Signal ---
		WB_ACK_O  <= WB_ACK_O_INT;

		--- Throttle ---
		WB_HALT_O <= '0'; -- yeay, we're at full speed!

		--- Error ---
		WB_ERR_O  <= '0'; -- nothing can go wrong ;)



end Behavioral;