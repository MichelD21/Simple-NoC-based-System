-- ######################################################
-- #          < STORM SoC by Stephan Nolting >          #
-- # ************************************************** #
-- #             Internal Memory Component              #
-- # ************************************************** #
-- # Last modified: 04.03.2012                          #
-- ######################################################

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;


entity MEMORY is
	generic	(
				MEM_SIZE      : natural := 256;  -- memory cells
				LOG2_MEM_SIZE : natural := 8;    -- log2(memory cells)
				OUTPUT_GATE   : boolean := FALSE -- output and-gate, might be necessary for some bus systems
			);
	port	(
				-- Wishbone Bus --
				WB_CLK_I      : in  STD_LOGIC; -- memory master clock
				WB_RST_I      : in  STD_LOGIC; -- high active sync reset
				WB_CTI_I      : in  STD_LOGIC_VECTOR(02 downto 0); -- cycle indentifier
				WB_TGC_I      : in  STD_LOGIC_VECTOR(06 downto 0); -- cycle tag
				WB_ADR_I      : in  STD_LOGIC_VECTOR(LOG2_MEM_SIZE-1 downto 0); -- adr in
				WB_DATA_I     : in  STD_LOGIC_VECTOR(31 downto 0); -- write data
				WB_DATA_O     : out STD_LOGIC_VECTOR(31 downto 0); -- read data
				WB_SEL_I      : in  STD_LOGIC_VECTOR(03 downto 0); -- data quantity
				WB_WE_I       : in  STD_LOGIC; -- write enable
				WB_STB_I      : in  STD_LOGIC; -- valid cycle
				WB_ACK_O      : out STD_LOGIC; -- acknowledge
				WB_HALT_O     : out STD_LOGIC; -- throttle master
				WB_ERR_O      : out STD_LOGIC  -- abnormal cycle termination
			);
end MEMORY;

architecture Behavioral of MEMORY is

	--- Buffer ---
	signal WB_ACK_O_INT : STD_LOGIC;
	signal WB_DATA_INT  : STD_LOGIC_VECTOR(31 downto 0);

	--- Memory Type ---
	type MEM_FILE_TYPE is array (0 to MEM_SIZE - 1) of STD_LOGIC_VECTOR(31 downto 0);

	--- INIT MEMORY IMAGE ---
	------------------------------------------------------
	signal MEM_FILE : MEM_FILE_TYPE :=
	(
		000000 => x"E10F1000",
000001 => x"E3C11080",
000002 => x"E121F001",
000003 => x"EB000000",
000004 => x"EAFFFFFE",
000005 => x"E3E01A01",
000006 => x"E3A02B01",
000007 => x"E5113FDB",
000008 => x"E5012FDF",
000009 => x"E5113FDB",
000010 => x"E3130B01",
000011 => x"E92D40F0",
000012 => x"1A000003",
000013 => x"E1A02001",
000014 => x"E5123FDB",
000015 => x"E3130B01",
000016 => x"0AFFFFFC",
000017 => x"E3A03C06",
000018 => x"E3A02B01",
000019 => x"E3E01A01",
000020 => x"E2833003",
000021 => x"E2822003",
000022 => x"E5013FDF",
000023 => x"E5012FDF",
000024 => x"E5113FDB",
000025 => x"E3130B01",
000026 => x"1A000003",
000027 => x"E1A02001",
000028 => x"E5123FDB",
000029 => x"E3130B01",
000030 => x"0AFFFFFC",
000031 => x"E3E01A01",
000032 => x"E3A03C06",
000033 => x"E3A02B01",
000034 => x"E5013FDF",
000035 => x"E5012FDF",
000036 => x"E5113FDB",
000037 => x"E3130B01",
000038 => x"1A000003",
000039 => x"E1A02001",
000040 => x"E5123FDB",
000041 => x"E3130B01",
000042 => x"0AFFFFFC",
000043 => x"E3E01A01",
000044 => x"E3A03C06",
000045 => x"E3A02B01",
000046 => x"E5013FDF",
000047 => x"E5012FDF",
000048 => x"E5113FDB",
000049 => x"E3130B01",
000050 => x"1A000003",
000051 => x"E1A02001",
000052 => x"E5123FDB",
000053 => x"E3130B01",
000054 => x"0AFFFFFC",
000055 => x"E3A03E63",
000056 => x"E3A02E43",
000057 => x"E3E01A01",
000058 => x"E2833002",
000059 => x"E2822002",
000060 => x"E5013FDF",
000061 => x"E5012FDF",
000062 => x"E5113FDB",
000063 => x"E3130B01",
000064 => x"1A000003",
000065 => x"E1A02001",
000066 => x"E5123FDB",
000067 => x"E3130B01",
000068 => x"0AFFFFFC",
000069 => x"E3A03E63",
000070 => x"E3A02E43",
000071 => x"E3E01A01",
000072 => x"E2833002",
000073 => x"E2822002",
000074 => x"E3A07000",
000075 => x"E5013FDF",
000076 => x"E59F6614",
000077 => x"E5012FDF",
000078 => x"E1A04007",
000079 => x"E3570031",
000080 => x"13A05000",
000081 => x"03A05001",
000082 => x"E3A01000",
000083 => x"E3E02A01",
000084 => x"E5123FDB",
000085 => x"E3510031",
000086 => x"13A00000",
000087 => x"02050001",
000088 => x"E3500000",
000089 => x"13A04001",
000090 => x"E3130B01",
000091 => x"E7D1E006",
000092 => x"1A000002",
000093 => x"E5123FDB",
000094 => x"E3130B01",
000095 => x"0AFFFFFC",
000096 => x"E1A0C404",
000097 => x"E38C3C06",
000098 => x"E183300E",
000099 => x"E3500000",
000100 => x"E1A03A83",
000101 => x"E1A03AA3",
000102 => x"E3E02A01",
000103 => x"13A00B01",
000104 => x"038C0B01",
000105 => x"E5023FDF",
000106 => x"E180300E",
000107 => x"13A04000",
000108 => x"E1A03A83",
000109 => x"E2811001",
000110 => x"11A0C004",
000111 => x"E1A03AA3",
000112 => x"E3E02A01",
000113 => x"E3510032",
000114 => x"E5023FDF",
000115 => x"1AFFFFDE",
000116 => x"E2877001",
000117 => x"E3570032",
000118 => x"E2866032",
000119 => x"1AFFFFD6",
000120 => x"E5123FDB",
000121 => x"E3130B01",
000122 => x"0AFFFFFC",
000123 => x"E38CCC06",
000124 => x"E38C3003",
000125 => x"E3802003",
000126 => x"E1A03A83",
000127 => x"E1A02A82",
000128 => x"E3E01A01",
000129 => x"E1A03AA3",
000130 => x"E1A02AA2",
000131 => x"E5013FDF",
000132 => x"E5012FDF",
000133 => x"E5113FDB",
000134 => x"E3130B01",
000135 => x"1A000003",
000136 => x"E1A02001",
000137 => x"E5123FDB",
000138 => x"E3130B01",
000139 => x"0AFFFFFC",
000140 => x"E38C3064",
000141 => x"E3802064",
000142 => x"E1A03A83",
000143 => x"E1A02A82",
000144 => x"E3E01A01",
000145 => x"E1A03AA3",
000146 => x"E1A02AA2",
000147 => x"E5013FDF",
000148 => x"E5012FDF",
000149 => x"E5113FDB",
000150 => x"E3130B01",
000151 => x"1A000003",
000152 => x"E1A02001",
000153 => x"E5123FDB",
000154 => x"E3130B01",
000155 => x"0AFFFFFC",
000156 => x"E1A03A8C",
000157 => x"E1A02A80",
000158 => x"E3E01A01",
000159 => x"E1A03AA3",
000160 => x"E1A02AA2",
000161 => x"E5013FDF",
000162 => x"E5012FDF",
000163 => x"E5113FDB",
000164 => x"E3130B01",
000165 => x"1A000003",
000166 => x"E1A02001",
000167 => x"E5123FDB",
000168 => x"E3130B01",
000169 => x"0AFFFFFC",
000170 => x"E3802032",
000171 => x"E38C3032",
000172 => x"E1A00A83",
000173 => x"E1A02A82",
000174 => x"E3E01A01",
000175 => x"E1A00AA0",
000176 => x"E1A02AA2",
000177 => x"E5010FDF",
000178 => x"E5012FDF",
000179 => x"E5113FDB",
000180 => x"E3130B01",
000181 => x"0AFFFFFC",
000182 => x"E3E03A01",
000183 => x"E5030FDF",
000184 => x"E59F6464",
000185 => x"E5032FDF",
000186 => x"E3A07000",
000187 => x"E3570031",
000188 => x"13A05000",
000189 => x"03A05001",
000190 => x"E3A01000",
000191 => x"E3E02A01",
000192 => x"E5123FDB",
000193 => x"E3510031",
000194 => x"13A00000",
000195 => x"02050001",
000196 => x"E3500000",
000197 => x"13A04001",
000198 => x"E3130B01",
000199 => x"E7D1E006",
000200 => x"1A000002",
000201 => x"E5123FDB",
000202 => x"E3130B01",
000203 => x"0AFFFFFC",
000204 => x"E1A0C404",
000205 => x"E38C3C06",
000206 => x"E183300E",
000207 => x"E3500000",
000208 => x"E1A03A83",
000209 => x"E1A03AA3",
000210 => x"E3E02A01",
000211 => x"13A00B01",
000212 => x"038C0B01",
000213 => x"E5023FDF",
000214 => x"E180300E",
000215 => x"13A0C000",
000216 => x"E1A03A83",
000217 => x"E2811001",
000218 => x"11A0400C",
000219 => x"E1A03AA3",
000220 => x"E3E02A01",
000221 => x"E3510032",
000222 => x"E5023FDF",
000223 => x"1AFFFFDE",
000224 => x"E2877001",
000225 => x"E3570032",
000226 => x"E2866032",
000227 => x"1AFFFFD6",
000228 => x"E5123FDB",
000229 => x"E3130B01",
000230 => x"0AFFFFFC",
000231 => x"E38C4C06",
000232 => x"E3843003",
000233 => x"E3802003",
000234 => x"E1A03A83",
000235 => x"E1A02A82",
000236 => x"E3E01A01",
000237 => x"E1A03AA3",
000238 => x"E1A02AA2",
000239 => x"E5013FDF",
000240 => x"E5012FDF",
000241 => x"E5113FDB",
000242 => x"E3130B01",
000243 => x"1A000003",
000244 => x"E1A02001",
000245 => x"E5123FDB",
000246 => x"E3130B01",
000247 => x"0AFFFFFC",
000248 => x"E3843064",
000249 => x"E3802064",
000250 => x"E1A03A83",
000251 => x"E1A02A82",
000252 => x"E3E01A01",
000253 => x"E1A03AA3",
000254 => x"E1A02AA2",
000255 => x"E5013FDF",
000256 => x"E5012FDF",
000257 => x"E5113FDB",
000258 => x"E3130B01",
000259 => x"1A000003",
000260 => x"E1A02001",
000261 => x"E5123FDB",
000262 => x"E3130B01",
000263 => x"0AFFFFFC",
000264 => x"E1A0EA84",
000265 => x"E1A0CA80",
000266 => x"E3E02A01",
000267 => x"E1A0EAAE",
000268 => x"E1A0CAAC",
000269 => x"E502EFDF",
000270 => x"E502CFDF",
000271 => x"E5123FDB",
000272 => x"E3130B01",
000273 => x"0AFFFFFC",
000274 => x"E3843032",
000275 => x"E3802032",
000276 => x"E1A03A83",
000277 => x"E1A02A82",
000278 => x"E3E01A01",
000279 => x"E1A03AA3",
000280 => x"E1A02AA2",
000281 => x"E5013FDF",
000282 => x"E5012FDF",
000283 => x"E5113FDB",
000284 => x"E3130B01",
000285 => x"1A000003",
000286 => x"E1A02001",
000287 => x"E5123FDB",
000288 => x"E3130B01",
000289 => x"0AFFFFFC",
000290 => x"E3E02A01",
000291 => x"E502EFDF",
000292 => x"E502CFDF",
000293 => x"E5123FDB",
000294 => x"E3130B01",
000295 => x"0AFFFFFC",
000296 => x"E3A03D1F",
000297 => x"E3A02D13",
000298 => x"E3E01A01",
000299 => x"E2833008",
000300 => x"E2822008",
000301 => x"E5013FDF",
000302 => x"E5012FDF",
000303 => x"E5113FDB",
000304 => x"E3130B01",
000305 => x"1A000003",
000306 => x"E1A02001",
000307 => x"E5123FDB",
000308 => x"E3130B01",
000309 => x"0AFFFFFC",
000310 => x"E3A03C06",
000311 => x"E3A02B01",
000312 => x"E3E01A01",
000313 => x"E2833003",
000314 => x"E2822003",
000315 => x"E5013FDF",
000316 => x"E5012FDF",
000317 => x"E5113FDB",
000318 => x"E3130B01",
000319 => x"1A000003",
000320 => x"E1A02001",
000321 => x"E5123FDB",
000322 => x"E3130B01",
000323 => x"0AFFFFFC",
000324 => x"E3A03D1B",
000325 => x"E3A02D13",
000326 => x"E3E01A01",
000327 => x"E2833008",
000328 => x"E2822008",
000329 => x"E5013FDF",
000330 => x"E5012FDF",
000331 => x"E5113FDB",
000332 => x"E3130B01",
000333 => x"1A000003",
000334 => x"E1A02001",
000335 => x"E5123FDB",
000336 => x"E3130B01",
000337 => x"0AFFFFFC",
000338 => x"E3A03D1B",
000339 => x"E3A02D13",
000340 => x"E3E01A01",
000341 => x"E2833008",
000342 => x"E2822008",
000343 => x"E5013FDF",
000344 => x"E5012FDF",
000345 => x"E5113FDB",
000346 => x"E3130B01",
000347 => x"1A000003",
000348 => x"E1A02001",
000349 => x"E5123FDB",
000350 => x"E3130B01",
000351 => x"0AFFFFFC",
000352 => x"E3E01A01",
000353 => x"E3A03C06",
000354 => x"E3A02B01",
000355 => x"E5013FDF",
000356 => x"E5012FDF",
000357 => x"E5113FDB",
000358 => x"E3130B01",
000359 => x"1A000003",
000360 => x"E1A02001",
000361 => x"E5123FDB",
000362 => x"E3130B01",
000363 => x"0AFFFFFC",
000364 => x"E3A03E63",
000365 => x"E3A02E43",
000366 => x"E3E01A01",
000367 => x"E2833002",
000368 => x"E2822002",
000369 => x"E5013FDF",
000370 => x"E5012FDF",
000371 => x"E5113FDB",
000372 => x"E3130B01",
000373 => x"1A000003",
000374 => x"E1A02001",
000375 => x"E5123FDB",
000376 => x"E3130B01",
000377 => x"0AFFFFFC",
000378 => x"E3A03E76",
000379 => x"E3A02E46",
000380 => x"E3E01A01",
000381 => x"E2833004",
000382 => x"E2822004",
000383 => x"E5013FDF",
000384 => x"E5012FDF",
000385 => x"E5113FDB",
000386 => x"E3130B01",
000387 => x"1A000003",
000388 => x"E1A02001",
000389 => x"E5123FDB",
000390 => x"E3130B01",
000391 => x"0AFFFFFC",
000392 => x"E3A03C06",
000393 => x"E3A02B01",
000394 => x"E3E01A01",
000395 => x"E2833003",
000396 => x"E2822003",
000397 => x"E5013FDF",
000398 => x"E5012FDF",
000399 => x"E5113FDB",
000400 => x"E3130B01",
000401 => x"1A000003",
000402 => x"E1A02001",
000403 => x"E5123FDB",
000404 => x"E3130B01",
000405 => x"0AFFFFFC",
000406 => x"E3A03E6D",
000407 => x"E3A02E4D",
000408 => x"E3E01A01",
000409 => x"E283300C",
000410 => x"E282200C",
000411 => x"E5013FDF",
000412 => x"E5012FDF",
000413 => x"E5113FDB",
000414 => x"E3130B01",
000415 => x"1A000003",
000416 => x"E1A02001",
000417 => x"E5123FDB",
000418 => x"E3130B01",
000419 => x"0AFFFFFC",
000420 => x"E3A03C06",
000421 => x"E3A02B01",
000422 => x"E3E01A01",
000423 => x"E283300A",
000424 => x"E282200A",
000425 => x"E5013FDF",
000426 => x"E5012FDF",
000427 => x"E5113FDB",
000428 => x"E3130B01",
000429 => x"1A000003",
000430 => x"E1A02001",
000431 => x"E5123FDB",
000432 => x"E3130B01",
000433 => x"0AFFFFFC",
000434 => x"E3E01A01",
000435 => x"E3A03C06",
000436 => x"E3A02B01",
000437 => x"E5013FDF",
000438 => x"E5012FDF",
000439 => x"E5113FDB",
000440 => x"E3130B01",
000441 => x"1A000003",
000442 => x"E1A02001",
000443 => x"E5123FDB",
000444 => x"E3130B01",
000445 => x"0AFFFFFC",
000446 => x"E3E01A01",
000447 => x"E3A03C06",
000448 => x"E3A02B01",
000449 => x"E5013FDF",
000450 => x"E5012FDF",
000451 => x"E5113FDB",
000452 => x"E3130B01",
000453 => x"1A000003",
000454 => x"E1A02001",
000455 => x"E5123FDB",
000456 => x"E3130B01",
000457 => x"0AFFFFFC",
000458 => x"E3A03E73",
000459 => x"E3A02E43",
000460 => x"E3E01A01",
000461 => x"E2833002",
000462 => x"E2822002",
000463 => x"E3A00000",
000464 => x"E5013FDF",
000465 => x"E5012FDF",
000466 => x"E8BD80F0",
000467 => x"00000850",
000468 => x"00000000",
000469 => x"00000000",
000470 => x"00000000",
000471 => x"00000000",
000472 => x"00000000",
000473 => x"00000000",
000474 => x"00000000",
000475 => x"00000000",
000476 => x"00000000",
000477 => x"00000000",
000478 => x"00000000",
000479 => x"00000000",
000480 => x"00000000",
000481 => x"00000000",
000482 => x"00000000",
000483 => x"00000000",
000484 => x"00000000",
000485 => x"00000000",
000486 => x"00000000",
000487 => x"00000000",
000488 => x"00000000",
000489 => x"00000000",
000490 => x"00000000",
000491 => x"00000000",
000492 => x"00000000",
000493 => x"00000000",
000494 => x"00000000",
000495 => x"00000000",
000496 => x"00000000",
000497 => x"00000000",
000498 => x"00000000",
000499 => x"00000000",
000500 => x"00000000",
000501 => x"00000000",
000502 => x"00000000",
000503 => x"00000000",
000504 => x"00000000",
000505 => x"00000000",
000506 => x"00000000",
000507 => x"00000000",
000508 => x"00000000",
000509 => x"00000000",
000510 => x"00000000",
000511 => x"00000000",
000512 => x"00000000",
000513 => x"00000000",
000514 => x"00000000",
000515 => x"00000000",
000516 => x"00000000",
000517 => x"00000000",
000518 => x"00000000",
000519 => x"00000000",
000520 => x"00000000",
000521 => x"00000000",
000522 => x"00000000",
000523 => x"00000000",
000524 => x"00000000",
000525 => x"00000000",
000526 => x"00000000",
000527 => x"00000000",
000528 => x"00000000",
000529 => x"00000000",
000530 => x"00000000",
000531 => x"00000000",
000532 => x"54540A00",
000533 => x"00000000",
000534 => x"00000A0A",
000535 => x"0A0A0000",
000536 => x"0A0A0A0B",
000537 => x"0B0B0B0B",
000538 => x"0B0A0A00",
000539 => x"0A0A0A0A",
000540 => x"0A0A0B4B",
000541 => x"0A000000",
000542 => x"00000000",
000543 => x"0000000A",
000544 => x"0A0B540C",
000545 => x"0A000000",
000546 => x"0A4C554D",
000547 => x"0A555554",
000548 => x"0A0A545C",
000549 => x"4C0B4C55",
000550 => x"55550C0B",
000551 => x"0A54540B",
000552 => x"0A0A0B0B",
000553 => x"5D540A00",
000554 => x"545C540A",
000555 => x"5C540000",
000556 => x"000A0A0C",
000557 => x"4B0B0A00",
000558 => x"00000B4D",
000559 => x"0B010B0B",
000560 => x"0B4C0A54",
000561 => x"4A0A4C0C",
000562 => x"0B0B4B0B",
000563 => x"55010B0B",
000564 => x"4B540A0A",
000565 => x"544C0B0A",
000566 => x"0B004C0A",
000567 => x"0A4D4A0B",
000568 => x"0000000A",
000569 => x"0A0C0A0A",
000570 => x"0A0A0000",
000571 => x"0A54F69D",
000572 => x"55FFF755",
000573 => x"004BF6F6",
000574 => x"0B559DF6",
000575 => x"F6F6074B",
000576 => x"0A07F654",
000577 => x"0A0B1455",
000578 => x"F607550A",
000579 => x"4CF6A54E",
000580 => x"F6070000",
000581 => x"00000A0B",
000582 => x"000A0A0A",
000583 => x"0A000A55",
000584 => x"F6AF4CFF",
000585 => x"A45E004B",
000586 => x"F6F60B55",
000587 => x"9DFFF6F6",
000588 => x"F60A0B07",
000589 => x"F6540A0B",
000590 => x"0C55F607",
000591 => x"9E0A4CFF",
000592 => x"A54EF6EE",
000593 => x"00000000",
000594 => x"0A0B000A",
000595 => x"4A0A0A00",
000596 => x"000AF6F6",
000597 => x"0AF60B01",
000598 => x"0A43F6F6",
000599 => x"4C559DF6",
000600 => x"A5F6FF9C",
000601 => x"0C07F654",
000602 => x"0A0B0D4D",
000603 => x"F6074C00",
000604 => x"4BFF9D56",
000605 => x"F6AE0000",
000606 => x"0000000A",
000607 => x"000A0A0A",
000608 => x"0A000A0A",
000609 => x"07FFFFF7",
000610 => x"0C0B0CAE",
000611 => x"F6F60754",
000612 => x"A5FFAE54",
000613 => x"F6AD4D08",
000614 => x"F6550A0C",
000615 => x"0D4BF6F6",
000616 => x"4B0C4BFF",
000617 => x"5C56FF08",
000618 => x"00000000",
000619 => x"0000000A",
000620 => x"0B0B0A00",
000621 => x"9D0AAEF6",
000622 => x"FF9C0B14",
000623 => x"0D07A4FF",
000624 => x"0755A5F6",
000625 => x"5C07F654",
000626 => x"0E08F655",
000627 => x"0A15565C",
000628 => x"F7F6544D",
000629 => x"4BFF5C56",
000630 => x"F6F70A00",
000631 => x"00000000",
000632 => x"000A0B4C",
000633 => x"0B0A5D53",
000634 => x"5DF6FF53",
000635 => x"0B150DF6",
000636 => x"5BFF0854",
000637 => x"9DF6EFF6",
000638 => x"F64B0E08",
000639 => x"F6550A55",
000640 => x"569DA5F6",
000641 => x"5C554CFF",
000642 => x"5C4EF6F7",
000643 => x"00000000",
000644 => x"00000A0B",
000645 => x"0C540C54",
000646 => x"00000BF6",
000647 => x"F64C0C15",
000648 => x"57084AF6",
000649 => x"085E9CFF",
000650 => x"08FF084C",
000651 => x"0EF6F655",
000652 => x"0A5D56F6",
000653 => x"9BF6AE56",
000654 => x"4CFF9D4D",
000655 => x"F6F70A0A",
000656 => x"0A0A0A00",
000657 => x"0A0B0C55",
000658 => x"0C0B0A00",
000659 => x"5DFFF60A",
000660 => x"0C5E1508",
000661 => x"0A08F654",
000662 => x"5CFF0808",
000663 => x"08530EF6",
000664 => x"F6550A56",
000665 => x"4CF653F6",
000666 => x"F7544CF6",
000667 => x"AE4EF6F7",
000668 => x"0A0A0A0A",
000669 => x"0A0A0C0C",
000670 => x"0C550C0B",
000671 => x"0A0AF6F6",
000672 => x"F69D0D15",
000673 => x"15F607F6",
000674 => x"F6AF5CF6",
000675 => x"9D0AF6F6",
000676 => x"5607FF56",
000677 => x"0B0C0BF6",
000678 => x"07F6080B",
000679 => x"01F65C57",
000680 => x"F6F70A0A",
000681 => x"0A0A0A0A",
000682 => x"0C0C0C55",
000683 => x"0C0B0A0A",
000684 => x"08F6F6A6",
000685 => x"0D1E15F6",
000686 => x"08FFF65E",
000687 => x"9DF69D0B",
000688 => x"F6F65608",
000689 => x"F6560B0C",
000690 => x"0AF608F6",
000691 => x"080B0CF6",
000692 => x"9D57F6F7",
000693 => x"0A0A0A0A",
000694 => x"0A0A155E",
000695 => x"5E0C0C0B",
000696 => x"0B55F6F6",
000697 => x"53F60C16",
000698 => x"55FF54F7",
000699 => x"FF5E5CFF",
000700 => x"F653F607",
000701 => x"5F07F64C",
000702 => x"54015DF6",
000703 => x"53F6F65C",
000704 => x"4CF6A456",
000705 => x"F6F70A0A",
000706 => x"0A0A0A0A",
000707 => x"151E550C",
000708 => x"0C0B0B15",
000709 => x"F6F654F6",
000710 => x"A7160DF6",
000711 => x"545CF656",
000712 => x"9DF6A507",
000713 => x"F6070D07",
000714 => x"F60A0A55",
000715 => x"A6F654F6",
000716 => x"F6A54DF6",
000717 => x"074CF6AD",
000718 => x"0A0A0A0A",
000719 => x"0A0A1455",
000720 => x"0D0C0C0B",
000721 => x"0C55F6A5",
000722 => x"5E08AE56",
000723 => x"EFF64D0B",
000724 => x"F65F5DF6",
000725 => x"F6F6F6B7",
000726 => x"AF07F6F6",
000727 => x"F656F6F6",
000728 => x"5607F6EE",
000729 => x"5508F6F6",
000730 => x"07530A0A",
000731 => x"0A0C0A0A",
000732 => x"0C675655",
000733 => x"5514554C",
000734 => x"074B5607",
000735 => x"EE015C08",
000736 => x"550B075E",
000737 => x"5DF608F6",
000738 => x"EF1CF608",
000739 => x"08080855",
000740 => x"9B0855A5",
000741 => x"08074D4B",
000742 => x"08084B54",
000743 => x"0B0B0B0B",
000744 => x"0A0A145E",
000745 => x"5E561515",
000746 => x"67550A0C",
000747 => x"160B0B0C",
000748 => x"0C0BA715",
000749 => x"0A56010B",
000750 => x"0A0A4C1E",
000751 => x"B70B0A5C",
000752 => x"0A560B0A",
000753 => x"4D0B0A0A",
000754 => x"0C540B0B",
000755 => x"540B0B0B",
000756 => x"0B0B0A0A",
000757 => x"0C155E5E",
000758 => x"1E676F6F",
000759 => x"67B71615",
000760 => x"15151516",
000761 => x"1515162F",
000762 => x"2F272727",
000763 => x"27272F1E",
000764 => x"1E1E1E15",
000765 => x"14151515",
000766 => x"15151515",
000767 => x"1455151E",
000768 => x"1514140C",
000769 => x"0B0A0C15",
000770 => x"5E5E1E67",
000771 => x"6F6F676F",
000772 => x"16151515",
000773 => x"15151515",
000774 => x"1E2F2F27",
000775 => x"6767272F",
000776 => x"2F1F1E1E",
000777 => x"1F151E15",
000778 => x"15151515",
000779 => x"16150C14",
000780 => x"151E1615",
000781 => x"150C0B0A",
000782 => x"1515151E",
000783 => x"1E676F6F",
000784 => x"271E1615",
000785 => x"15151515",
000786 => x"16161E6F",
000787 => x"2F2F6F6F",
000788 => x"6F6F6F6F",
000789 => x"B766671E",
000790 => x"6F6F1E15",
000791 => x"151E5F16",
000792 => x"15151515",
000793 => x"150C140C",
000794 => x"0B0A1515",
000795 => x"151E1E27",
000796 => x"6F6F1E1E",
000797 => x"16151515",
000798 => x"15161E1E",
000799 => x"1F6F2F6F",
000800 => x"6FB7B76F",
000801 => x"6FAFB7B7",
000802 => x"B71E2727",
000803 => x"6715151E",
000804 => x"1F161515",
000805 => x"15151555",
000806 => x"14140B0A",
000807 => x"1515551E",
000808 => x"1F1F6F6F",
000809 => x"1F1F1E15",
000810 => x"1515151E",
000811 => x"1E1E272F",
000812 => x"77BFEF5D",
000813 => x"EEF6F6B6",
000814 => x"AFAEF66F",
000815 => x"272F6F1E",
000816 => x"1E1E6F27",
000817 => x"1E165656",
000818 => x"0E564D15",
000819 => x"0C0A1515",
000820 => x"551E1F1F",
000821 => x"6F6F1F1F",
000822 => x"1E151515",
000823 => x"151E1E1E",
000824 => x"272F77BF",
000825 => x"EF5DEEF6",
000826 => x"F6B6AFAE",
000827 => x"F66F272F",
000828 => x"6F1E1E1E",
000829 => x"6F271E16",
000830 => x"56560E56",
000831 => x"4D150C0A",
000832 => x"150C0D16",
000833 => x"161F2F6F",
000834 => x"1F1F1E16",
000835 => x"161E1F1F",
000836 => x"2727276F",
000837 => x"6FF6F65C",
000838 => x"07EFB7B7",
000839 => x"A5F6F6B7",
000840 => x"6F6F6F27",
000841 => x"272F7727",
000842 => x"1F1E0E4E",
000843 => x"4E4D4E15",
000844 => x"0C0B1555",
000845 => x"4D56561E",
000846 => x"2F2F2727",
000847 => x"271E1E1F",
000848 => x"1F272727",
000849 => x"2F776FF6",
000850 => x"F608F6AF",
000851 => x"67AFF6F6",
000852 => x"F6AF6F6F",
000853 => x"6F6F2F6F",
000854 => x"77271E1F",
000855 => x"0E0E0E4E",
000856 => x"5515140C",
000857 => x"154D4E4E",
000858 => x"4E5E2F2F",
000859 => x"271F2727",
000860 => x"271E2727",
000861 => x"27272F6F",
000862 => x"66F6F6F6",
000863 => x"B7675F67",
000864 => x"EFF6F6AF",
000865 => x"67672F77",
000866 => x"6F777727",
000867 => x"1E1F0E4E",
000868 => x"0E0D1515",
000869 => x"140C1E0D",
000870 => x"4D4D4D56",
000871 => x"2F272727",
000872 => x"27272727",
000873 => x"27272727",
000874 => x"2767555D",
000875 => x"A55D551F",
000876 => x"1F5F56AF",
000877 => x"EF55561E",
000878 => x"77777777",
000879 => x"7727275F",
000880 => x"0D0D0D15",
000881 => x"67151415",
000882 => x"1E0D4D4D",
000883 => x"4D152727",
000884 => x"27272727",
000885 => x"27672727",
000886 => x"2727275E",
000887 => x"1554544C",
000888 => x"0D1F1F5F",
000889 => x"55A6AF55",
000890 => x"56167777",
000891 => x"77777727",
000892 => x"675F0D0D",
000893 => x"0D155E15",
000894 => x"141D1E56",
000895 => x"550D0D56",
000896 => x"671F2727",
000897 => x"6F6F2767",
000898 => x"27272727",
000899 => x"670D0D01",
000900 => x"0C010117",
000901 => x"17570E0C",
000902 => x"4D0D0D56",
000903 => x"6F777777",
000904 => x"772F671E",
000905 => x"014D151E",
000906 => x"5E14141E",
000907 => x"275E560D",
000908 => x"4D0D155F",
000909 => x"2727776F",
000910 => x"2F2F272F",
000911 => x"27675F4D",
000912 => x"0C010C0C",
000913 => x"010D570E",
000914 => x"0C0B0C0C",
000915 => x"0C4D1F77",
000916 => x"2F2F2F67",
000917 => x"1E0D0D0D",
000918 => x"5E1E1515",
000919 => x"141E275E",
000920 => x"560D4D0D",
000921 => x"155F2727",
000922 => x"776F2F2F",
000923 => x"272F2767",
000924 => x"5F4D0C01",
000925 => x"0C0C010D",
000926 => x"570E0C0B",
000927 => x"0C0C0C4D",
000928 => x"1F772F2F",
000929 => x"2F671E0D",
000930 => x"0D0D5E1E",
000931 => x"1515141E",
000932 => x"27272F6F",
000933 => x"67550D0D",
000934 => x"67672F2F",
000935 => x"2F2F6F1E",
000936 => x"56564E0C",
000937 => x"0B0B0B0B",
000938 => x"0B0B0B0A",
000939 => x"0A0A0A0A",
000940 => x"0B0C4E56",
000941 => x"1F6F6715",
000942 => x"0D0D155E",
000943 => x"1E676715",
000944 => x"1E67272F",
000945 => x"2F6F6F15",
000946 => x"4E0D5E77",
000947 => x"2F2F2F2F",
000948 => x"6F56564E",
000949 => x"4E0C0B0C",
000950 => x"0C0C4C4C",
000951 => x"4C0B0B0B",
000952 => x"0B0A0B0C",
000953 => x"4E571F6F",
000954 => x"270D4D0D",
000955 => x"165E1E27",
000956 => x"1655151E",
000957 => x"2F2F2F77",
000958 => x"77670D4D",
000959 => x"0D1E676F",
000960 => x"2F376F16",
000961 => x"0E0E4E0C",
000962 => x"0D0C0D0D",
000963 => x"0C0D0D0D",
000964 => x"0D0D0C0C",
000965 => x"0C0D4E56",
000966 => x"5F6F164D",
000967 => x"4D0D5E1E",
000968 => x"1E151515",
000969 => x"15152F2F",
000970 => x"3777776F",
000971 => x"0D4D0D15",
000972 => x"672F2F37",
000973 => x"6F5F0E0E",
000974 => x"4E0C0D0C",
000975 => x"0D0D0D0D",
000976 => x"0D0D0D0D",
000977 => x"0D0C0C0D",
000978 => x"4E565E67",
000979 => x"164D4D0D",
000980 => x"671E1515",
000981 => x"0D151515",
000982 => x"37373737",
000983 => x"37775F16",
000984 => x"4D0D1577",
000985 => x"77777767",
000986 => x"0D0D0D01",
000987 => x"0101010C",
000988 => x"0C0C0C01",
000989 => x"0D0D0D0D",
000990 => x"0D4D4D0D",
000991 => x"4E564E0D",
000992 => x"0D5E1E1E",
000993 => x"160C0C15",
000994 => x"15153737",
000995 => x"37373737",
000996 => x"671E560D",
000997 => x"0D6F7777",
000998 => x"77670D0D",
000999 => x"0D010101",
001000 => x"010C0101",
001001 => x"0C010D01",
001002 => x"0D0D0D0D",
001003 => x"4D4D0D4E",
001004 => x"4E0D565F",
001005 => x"1E15150C",
001006 => x"0C0C1515",
001007 => x"3777372F",
001008 => x"2F2F776F",
001009 => x"160E4D0D",
001010 => x"6F6F2F6F",
001011 => x"5E4C0C0D",
001012 => x"010C0C01",
001013 => x"01010C0D",
001014 => x"0D0D4D0D",
001015 => x"0C01014D",
001016 => x"4D4E0D16",
001017 => x"67271516",
001018 => x"150C0B0C",
001019 => x"67273737",
001020 => x"7737372F",
001021 => x"3777160E",
001022 => x"0D0D1527",
001023 => x"2F6F670C",
001024 => x"0C4D010C",
001025 => x"0C01010C",
001026 => x"0C0D0D0D",
001027 => x"0D0C0101",
001028 => x"0C0D0D4E",
001029 => x"0D676727",
001030 => x"151E150C",
001031 => x"0C0C6767",
001032 => x"3F7F7737",
001033 => x"372F3777",
001034 => x"5F560D4D",
001035 => x"0D15272F",
001036 => x"670C0101",
001037 => x"010C0C01",
001038 => x"010C0C0D",
001039 => x"0D0D0D01",
001040 => x"010C4C0D",
001041 => x"0D0D566F",
001042 => x"2F271E15",
001043 => x"1E150C55",
001044 => x"6727FB7F",
001045 => x"772F2F27",
001046 => x"2F376F5E",
001047 => x"164D0D0E",
001048 => x"1F6F670C",
001049 => x"0D4D0C0C",
001050 => x"0C010C01",
001051 => x"010D4D0D",
001052 => x"0D010C0C",
001053 => x"0C0D0D0D",
001054 => x"1E6F2F6F",
001055 => x"1F1E165E",
001056 => x"155E6F6F",
001057 => x"3F7F7737",
001058 => x"2F2F2F2F",
001059 => x"6F67164D",
001060 => x"4D0D166F",
001061 => x"670C0D4D",
001062 => x"0C0C0C0C",
001063 => x"0C0C010D",
001064 => x"4D0D0D01",
001065 => x"0C010C0D",
001066 => x"4D0D1E2F",
001067 => x"2F6F1E1F",
001068 => x"155E1567",
001069 => x"6F6FFBFB",
001070 => x"7F777F2F",
001071 => x"372F7F7F",
001072 => x"77564E4E",
001073 => x"0D0C0D4D",
001074 => x"0C4D0D0C",
001075 => x"0D4D0C01",
001076 => x"0C0D0C01",
001077 => x"0C0C0C01",
001078 => x"4C4D0D15",
001079 => x"7737772F",
001080 => x"271E2716",
001081 => x"16672777",
001082 => x"FBFB7F77",
001083 => x"7F2F372F",
001084 => x"7F7F7756",
001085 => x"4E4E0D0C",
001086 => x"0D4D0C4D",
001087 => x"0D0C0D4D",
001088 => x"0C010C0D",
001089 => x"0C010C0C",
001090 => x"0C014C4D",
001091 => x"0D157737",
001092 => x"772F271E",
001093 => x"27161667",
001094 => x"27773F37",
001095 => x"2F27275F",
001096 => x"27277F7F",
001097 => x"7F771E56",
001098 => x"150D0C01",
001099 => x"0C0C0C01",
001100 => x"0101010C",
001101 => x"010C0101",
001102 => x"010C0C01",
001103 => x"0C561E77",
001104 => x"77772F2F",
001105 => x"27675E15",
001106 => x"15151F67",
001107 => x"37372F27",
001108 => x"271E2727",
001109 => x"7F7F7F77",
001110 => x"2656160D",
001111 => x"0C010C01",
001112 => x"0C010C01",
001113 => x"010C0101",
001114 => x"010C0C0D",
001115 => x"0D0C0D56",
001116 => x"1E777777",
001117 => x"2F2F2727",
001118 => x"6715150D",
001119 => x"1E67372F",
001120 => x"2F2F2716",
001121 => x"1E277F7F",
001122 => x"3F777767",
001123 => x"160D0C01",
001124 => x"010C4C0C",
001125 => x"0C0C010C",
001126 => x"0101010C",
001127 => x"010D0D0D",
001128 => x"0D556777",
001129 => x"772F6F6F",
001130 => x"671E675E",
001131 => x"AF0C1567",
001132 => x"372F2727",
001133 => x"271E1F27",
001134 => x"77373777",
001135 => x"7F771E0D",
001136 => x"0C0C0C0C",
001137 => x"0C0C4D0C",
001138 => x"010C0101",
001139 => x"0C0D0D4E",
001140 => x"4D014D0D",
001141 => x"77772F27",
001142 => x"2727671F",
001143 => x"6F5F550C",
001144 => x"0C15376F",
001145 => x"2727271E",
001146 => x"1F677777",
001147 => x"777F7F77",
001148 => x"665F4D4C",
001149 => x"4C0D0C4D",
001150 => x"4D0D0D0D",
001151 => x"0C0C0C0C",
001152 => x"0D0D550D",
001153 => x"555E6F77",
001154 => x"6F27676F",
001155 => x"67676767",
001156 => x"150B0C14",
others => x"F0013007"

);
	------------------------------------------------------

begin

	-- STORM data/instruction memory -----------------------------------------------------------------------
	-- --------------------------------------------------------------------------------------------------------
		MEM_FILE_ACCESS: process(WB_CLK_I)
		begin
			--- Sync Write ---
			if rising_edge(WB_CLK_I) then

				--- Data Read/Write ---
				if (WB_STB_I = '1') then
					if (WB_WE_I = '1') then
						MEM_FILE(to_integer(unsigned(WB_ADR_I))) <= WB_DATA_I;
					end if;
					WB_DATA_INT <= MEM_FILE(to_integer(unsigned(WB_ADR_I)));
				end if;

				--- ACK Control ---
				if (WB_RST_I = '1') then
					WB_ACK_O_INT <= '0';
				elsif (WB_CTI_I = "000") or (WB_CTI_I = "111") then
					WB_ACK_O_INT <= WB_STB_I and (not WB_ACK_O_INT);
				else
					WB_ACK_O_INT <= WB_STB_I;
				end if;

			end if;
		end process MEM_FILE_ACCESS;

		--- Output Gate ---
		WB_DATA_O <= WB_DATA_INT when (OUTPUT_GATE = FALSE) or ((OUTPUT_GATE = TRUE) and (WB_STB_I = '1')) else (others => '0');

		--- ACK Signal ---
		WB_ACK_O  <= WB_ACK_O_INT;

		--- Throttle ---
		WB_HALT_O <= '0'; -- yeay, we're at full speed!

		--- Error ---
		WB_ERR_O  <= '0'; -- nothing can go wrong ;)



end Behavioral;