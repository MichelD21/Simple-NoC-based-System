-- ######################################################
-- #          < STORM SoC by Stephan Nolting >          #
-- # ************************************************** #
-- #             Internal Memory Component              #
-- # ************************************************** #
-- # Last modified: 04.03.2012                          #
-- ######################################################

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;


entity MEMORY is
	generic	(
				MEM_SIZE      : natural := 256;  -- memory cells
				LOG2_MEM_SIZE : natural := 8;    -- log2(memory cells)
				OUTPUT_GATE   : boolean := FALSE -- output and-gate, might be necessary for some bus systems
			);
	port	(
				-- Wishbone Bus --
				WB_CLK_I      : in  STD_LOGIC; -- memory master clock
				WB_RST_I      : in  STD_LOGIC; -- high active sync reset
				WB_CTI_I      : in  STD_LOGIC_VECTOR(02 downto 0); -- cycle indentifier
				WB_TGC_I      : in  STD_LOGIC_VECTOR(06 downto 0); -- cycle tag
				WB_ADR_I      : in  STD_LOGIC_VECTOR(LOG2_MEM_SIZE-1 downto 0); -- adr in
				WB_DATA_I     : in  STD_LOGIC_VECTOR(31 downto 0); -- write data
				WB_DATA_O     : out STD_LOGIC_VECTOR(31 downto 0); -- read data
				WB_SEL_I      : in  STD_LOGIC_VECTOR(03 downto 0); -- data quantity
				WB_WE_I       : in  STD_LOGIC; -- write enable
				WB_STB_I      : in  STD_LOGIC; -- valid cycle
				WB_ACK_O      : out STD_LOGIC; -- acknowledge
				WB_HALT_O     : out STD_LOGIC; -- throttle master
				WB_ERR_O      : out STD_LOGIC  -- abnormal cycle termination
			);
end MEMORY;

architecture Behavioral of MEMORY is

	--- Buffer ---
	signal WB_ACK_O_INT : STD_LOGIC;
	signal WB_DATA_INT  : STD_LOGIC_VECTOR(31 downto 0);

	--- Memory Type ---
	type MEM_FILE_TYPE is array (0 to MEM_SIZE - 1) of STD_LOGIC_VECTOR(31 downto 0);

	--- INIT MEMORY IMAGE ---
	------------------------------------------------------
	signal MEM_FILE : MEM_FILE_TYPE :=
	(
		000000 => x"E10F1000",
000001 => x"E3C11080",
000002 => x"E121F001",
000003 => x"EB000000",
000004 => x"EAFFFFFE",
000005 => x"E3E03A01",
000006 => x"E5132FDB",
000007 => x"E3A02B01",
000008 => x"E92D40F0",
000009 => x"E5032FDF",
000010 => x"E59F7108",
000011 => x"E3A06000",
000012 => x"E087E286",
000013 => x"E3A0C000",
000014 => x"E3865C06",
000015 => x"E3864B01",
000016 => x"E3E02A01",
000017 => x"E5123FDB",
000018 => x"E3130B01",
000019 => x"0AFFFFFC",
000020 => x"E3A03C06",
000021 => x"E3A02B01",
000022 => x"E3E01A01",
000023 => x"E2833003",
000024 => x"E2822003",
000025 => x"E5013FDF",
000026 => x"E5012FDF",
000027 => x"E5113FDB",
000028 => x"E3130B01",
000029 => x"1A000003",
000030 => x"E1A02001",
000031 => x"E5123FDB",
000032 => x"E3130B01",
000033 => x"0AFFFFFC",
000034 => x"E1A03A85",
000035 => x"E1A02A84",
000036 => x"E3E01A01",
000037 => x"E1A03AA3",
000038 => x"E1A02AA2",
000039 => x"E5013FDF",
000040 => x"E5012FDF",
000041 => x"E5113FDB",
000042 => x"E3130B01",
000043 => x"1A000003",
000044 => x"E1A02001",
000045 => x"E5123FDB",
000046 => x"E3130B01",
000047 => x"0AFFFFFC",
000048 => x"E38C3C06",
000049 => x"E38C2B01",
000050 => x"E1A03A83",
000051 => x"E1A02A82",
000052 => x"E3E01A01",
000053 => x"E1A03AA3",
000054 => x"E1A02AA2",
000055 => x"E5013FDF",
000056 => x"E5012FDF",
000057 => x"E5113FDB",
000058 => x"E3130B01",
000059 => x"E5DE0000",
000060 => x"1A000003",
000061 => x"E1A02001",
000062 => x"E5123FDB",
000063 => x"E3130B01",
000064 => x"0AFFFFFC",
000065 => x"E28CC001",
000066 => x"E3E02A01",
000067 => x"E3801B01",
000068 => x"E3803C07",
000069 => x"E35C0020",
000070 => x"E5023FDF",
000071 => x"E28EE001",
000072 => x"E5021FDF",
000073 => x"1AFFFFC5",
000074 => x"E2866001",
000075 => x"E3560018",
000076 => x"1AFFFFBE",
000077 => x"EAFFFFFE",
000078 => x"0000023C",
000079 => x"00000000",
000080 => x"00000000",
000081 => x"00000000",
000082 => x"00000000",
000083 => x"00000000",
000084 => x"00000000",
000085 => x"00000000",
000086 => x"00000000",
000087 => x"00000000",
000088 => x"00000000",
000089 => x"00000000",
000090 => x"00000000",
000091 => x"00000000",
000092 => x"00000000",
000093 => x"00000000",
000094 => x"00000000",
000095 => x"00000000",
000096 => x"00000000",
000097 => x"00000000",
000098 => x"00000000",
000099 => x"00000000",
000100 => x"00000000",
000101 => x"00000000",
000102 => x"00000000",
000103 => x"00000000",
000104 => x"00000000",
000105 => x"00000000",
000106 => x"00000000",
000107 => x"00000000",
000108 => x"00000000",
000109 => x"00000000",
000110 => x"00000000",
000111 => x"00000000",
000112 => x"00000000",
000113 => x"00000000",
000114 => x"00000000",
000115 => x"00000000",
000116 => x"00000000",
000117 => x"00000000",
000118 => x"00000000",
000119 => x"00000000",
000120 => x"00000000",
000121 => x"00000000",
000122 => x"00000000",
000123 => x"00000000",
000124 => x"00000000",
000125 => x"00000000",
000126 => x"00000000",
000127 => x"00000000",
000128 => x"00000000",
000129 => x"00000000",
000130 => x"00000000",
000131 => x"00000000",
000132 => x"00000000",
000133 => x"00000000",
000134 => x"00000000",
000135 => x"00000000",
000136 => x"00000000",
000137 => x"00000000",
000138 => x"00000000",
000139 => x"00000000",
000140 => x"00000000",
000141 => x"00000000",
000142 => x"00000000",
000143 => x"0909ECEC",
000144 => x"ECECECF4",
000145 => x"F5F5F5F5",
000146 => x"090909F6",
000147 => x"F6090909",
000148 => x"09070909",
000149 => x"F6F6F6F6",
000150 => x"F6090909",
000151 => x"09090909",
000152 => x"ECECECF4",
000153 => x"ECECECF5",
000154 => x"F4F509A4",
000155 => x"A4090909",
000156 => x"09090909",
000157 => x"09090909",
000158 => x"09090909",
000159 => x"F5090909",
000160 => x"F5F5F5F5",
000161 => x"F4F4F5EC",
000162 => x"ECEC9241",
000163 => x"00A4EDF4",
000164 => x"F4090909",
000165 => x"09090909",
000166 => x"09090909",
000167 => x"09090909",
000168 => x"09090909",
000169 => x"09F40909",
000170 => x"09095200",
000171 => x"00F7EDEC",
000172 => x"E3ECECEC",
000173 => x"ECECECED",
000174 => x"09090909",
000175 => x"09090909",
000176 => x"09090909",
000177 => x"F5F5F509",
000178 => x"09090949",
000179 => x"51090909",
000180 => x"090909F4",
000181 => x"ECECE3A3",
000182 => x"E3E3E4EC",
000183 => x"F5F509F5",
000184 => x"09090909",
000185 => x"090909EC",
000186 => x"E4EC0909",
000187 => x"EC090909",
000188 => x"09090909",
000189 => x"0909F5F5",
000190 => x"ECECECEC",
000191 => x"09090909",
000192 => x"09F5F5F5",
000193 => x"F50909DA",
000194 => x"919189EC",
000195 => x"ECECEBEC",
000196 => x"ECF509F4",
000197 => x"F5090909",
000198 => x"09ECECEC",
000199 => x"09090909",
000200 => x"09090909",
000201 => x"F5ECE2DA",
000202 => x"914040DA",
000203 => x"9BF5F4EB",
000204 => x"F4ECECEC",
000205 => x"EC090909",
000206 => x"09F5ECEC",
000207 => x"F5F50909",
000208 => x"0909F4EC",
000209 => x"EDE3DAE3",
000210 => x"91480049",
000211 => x"EC09F409",
000212 => x"07F50909",
000213 => x"ECECECEC",
000214 => x"ECECEC09",
000215 => x"F5F5EDED",
000216 => x"F5F5ECEC",
000217 => x"EC484849",
000218 => x"4800A392",
000219 => x"92ECEBA3",
000220 => x"A3E3F4EC",
000221 => x"ECECECEC",
000222 => x"E3E3E3E3",
000223 => x"F5EDECEC",
000224 => x"ECEDEDED",
000225 => x"ED000000",
000226 => x"0000ED09",
000227 => x"899A0909",
000228 => x"ECE3E3EC",
000229 => x"E3E3ECEC",
000230 => x"ECECF5F4",
000231 => x"0909F5F5",
000232 => x"EDEDECEC",
000233 => x"ED490000",
000234 => x"000000ED",
000235 => x"0992A209",
000236 => x"09F50909",
000237 => x"ECE4ECEC",
000238 => x"E3E3ECEC",
000239 => x"09090909",
000240 => x"09090909",
000241 => x"09ED0000",
000242 => x"00000049",
000243 => x"EDF59B4A",
000244 => x"E507EDEC",
000245 => x"F5ECEDF5",
000246 => x"ECECECF5",
000247 => x"09090909",
000248 => x"09090909",
000249 => x"09F6A400",
000250 => x"00520000",
000251 => x"49F5F552",
000252 => x"52EE09F5",
000253 => x"F5EDECEC",
000254 => x"ECECEDF5",
000255 => x"F6F60909",
000256 => x"09090909",
000257 => x"0909A300",
000258 => x"9BF6F500",
000259 => x"49F50907",
000260 => x"EDEDF5ED",
000261 => x"EDECECEC",
000262 => x"ECECECEC",
000263 => x"FFFFF609",
000264 => x"0909F5F5",
000265 => x"09AC0052",
000266 => x"F6090949",
000267 => x"00090909",
000268 => x"0909F509",
000269 => x"F5ECEDED",
000270 => x"EDECEDF5",
000271 => x"0909FFFF",
000272 => x"FFF60907",
000273 => x"074900E4",
000274 => x"09090951",
000275 => x"00ED0909",
000276 => x"07F50909",
000277 => x"09090909",
000278 => x"F5F5ECEC",
000279 => x"A3E3ED09",
000280 => x"F6F6F6FF",
000281 => x"ED92EDED",
000282 => x"A3E3E39A",
000283 => x"00AC0909",
000284 => x"09090909",
000285 => x"09090909",
000286 => x"09090909",
000287 => x"ECE39BA3",
000288 => x"A3E3E3E4",
000289 => x"E4ECFFFF",
000290 => x"0809ED9B",
000291 => x"0092ECEC",
000292 => x"ECECE3EC",
000293 => x"F5F50909",
000294 => x"09090909",
000295 => x"0909EDED",
000296 => x"ECE39A91",
000297 => x"49529CF7",
000298 => x"08F6FF07",
000299 => x"000048A3",
000300 => x"ECA3DBDA",
000301 => x"E3E3EBEB",
000302 => x"ECF5F4F5",
000303 => x"09090909",
000304 => x"09F5F5F5",
000305 => x"51004952",
000306 => x"929BA4A4",
000307 => x"525353B7",
000308 => x"BFB70807",
000309 => x"07F7EDF7",
000310 => x"E4E4E3E3",
000311 => x"09090909",
000312 => x"09090909",
000313 => x"9A4091EC",
000314 => x"ECE3A300",
000315 => x"4952A5AF",
000316 => x"6E6FB7BF",
000317 => x"B7B7BFB7",
000318 => x"07F7E3E3",
000319 => x"09090909",
000320 => x"09090909",
000321 => x"9A48A3EC",
000322 => x"F409A300",
000323 => x"E3E4E4EC",
000324 => x"A49B9B9A",
000325 => x"E39B9B9B",
000326 => x"DBE3E3EC",
000327 => x"09090909",
000328 => x"090909EC",
000329 => x"9249A4ED",
000330 => x"F5EC5152",
000331 => x"F5F50909",
000332 => x"090709F5",
000333 => x"ECECE4EC",
000334 => x"ECECECE3",
others => x"F0013007"


);
	------------------------------------------------------

begin

	-- STORM data/instruction memory -----------------------------------------------------------------------
	-- --------------------------------------------------------------------------------------------------------
		MEM_FILE_ACCESS: process(WB_CLK_I)
		begin
			--- Sync Write ---
			if rising_edge(WB_CLK_I) then

				--- Data Read/Write ---
				if (WB_STB_I = '1') then
					if (WB_WE_I = '1') then
						MEM_FILE(to_integer(unsigned(WB_ADR_I))) <= WB_DATA_I;
					end if;
					WB_DATA_INT <= MEM_FILE(to_integer(unsigned(WB_ADR_I)));
				end if;

				--- ACK Control ---
				if (WB_RST_I = '1') then
					WB_ACK_O_INT <= '0';
				elsif (WB_CTI_I = "000") or (WB_CTI_I = "111") then
					WB_ACK_O_INT <= WB_STB_I and (not WB_ACK_O_INT);
				else
					WB_ACK_O_INT <= WB_STB_I;
				end if;

			end if;
		end process MEM_FILE_ACCESS;

		--- Output Gate ---
		WB_DATA_O <= WB_DATA_INT when (OUTPUT_GATE = FALSE) or ((OUTPUT_GATE = TRUE) and (WB_STB_I = '1')) else (others => '0');

		--- ACK Signal ---
		WB_ACK_O  <= WB_ACK_O_INT;

		--- Throttle ---
		WB_HALT_O <= '0'; -- yeay, we're at full speed!

		--- Error ---
		WB_ERR_O  <= '0'; -- nothing can go wrong ;)



end Behavioral;